
module FA_513 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_693 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_692 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_691 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_690 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_689 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_688 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_687 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_686 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_685 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_684 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_683 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_682 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_681 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_680 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_679 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_678 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_677 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_676 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_675 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_674 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_673 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_672 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_671 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_670 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_669 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_668 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_667 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_666 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_665 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_664 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_663 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_662 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_661 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_660 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_659 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_658 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_657 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_656 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_655 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_654 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_653 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_652 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_651 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_650 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_649 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_648 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_647 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_646 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_645 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_644 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_643 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_642 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_641 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_640 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_639 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_638 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_637 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_635 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_634 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_633 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_631 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_630 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_629 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_628 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_627 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_626 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_625 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_624 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_623 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_622 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_621 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_620 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_619 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_618 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_617 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_616 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_615 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_614 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_613 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_612 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_611 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_610 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_609 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_608 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_607 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_606 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_605 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_604 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_603 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_602 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_601 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_600 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_599 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_598 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_597 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_596 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_595 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_594 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_593 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_592 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_591 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_590 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_589 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_588 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_587 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_586 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_585 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_584 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_583 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_582 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_581 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_580 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_579 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_578 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_577 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_576 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_575 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_574 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_573 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_572 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_569 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_568 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_561 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_557 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_550 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_548 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_545 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_542 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_534 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_533 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_532 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_530 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_529 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_528 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_526 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_521 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_518 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_517 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module FA_514 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
  INV_X1 U2 ( .A(n18), .ZN(Co) );
endmodule


module FA_512 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n18, n19;

  XOR2_X1 U3 ( .A(Ci), .B(n19), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n19) );
  INV_X1 U1 ( .A(n18), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n19), .B2(Ci), .ZN(n18) );
endmodule


module PG_97 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_96 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_92 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_91 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_90 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_89 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_88 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_87 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_80 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_79 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_78 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_77 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_76 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_74 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_73 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_70 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_69 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_65 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_64 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_63 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_62 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_61 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_60 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_58 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_41 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_40 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_85 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_84 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_83 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_81 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_75 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_72 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_71 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_68 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_67 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_66 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_59 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_57 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_56 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module PG_30 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_28 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n10;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n10) );
endmodule


module G_26 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n10) );
endmodule


module G_25 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n10) );
endmodule


module G_24 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n10) );
endmodule


module G_23 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n10) );
endmodule


module G_22 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n10) );
endmodule


module G_21 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n10) );
endmodule


module G_20 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n10) );
endmodule


module G_19 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n10) );
endmodule


module G_10 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n10;

  INV_X1 U1 ( .A(n10), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n10) );
endmodule


module PGblock_120 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_119 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_118 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_117 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_116 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_115 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_114 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_113 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_112 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_111 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_110 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_109 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_108 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_107 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_106 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_105 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_104 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_103 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_102 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_101 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_100 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_99 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_98 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_97 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_96 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_95 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_94 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_93 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_92 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_91 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_90 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_89 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_88 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_87 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_86 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_85 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_84 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_83 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_82 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_81 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_80 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_79 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_78 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_77 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_76 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_75 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_74 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_73 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_72 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_71 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_70 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_69 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_68 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_67 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_66 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_65 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_62 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_60 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_59 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_58 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_54 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_52 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_50 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_48 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_47 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_46 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_45 ( A, B, G, P );
  input A, B;
  output G, P;
  wire   n1;

  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  CLKBUF_X1 U1 ( .A(B), .Z(n1) );
  AND2_X1 U3 ( .A1(n1), .A2(A), .ZN(G) );
endmodule


module PGblock_44 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_43 ( A, B, G, P );
  input A, B;
  output G, P;
  wire   n1;

  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  CLKBUF_X1 U1 ( .A(B), .Z(n1) );
  AND2_X1 U3 ( .A1(n1), .A2(A), .ZN(G) );
endmodule


module PGblock_42 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_41 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_40 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_39 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_38 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_37 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_36 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_35 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_34 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_33 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module RegEn_Nbit32_2 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;


  FD_EN_69 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_68 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_67 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_66 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_65 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
  FD_EN_64 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[5]) );
  FD_EN_63 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[6]) );
  FD_EN_62 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[7]) );
  FD_EN_61 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[8]) );
  FD_EN_60 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[9]) );
  FD_EN_59 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[10]) );
  FD_EN_58 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[11]) );
  FD_EN_57 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[12]) );
  FD_EN_56 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[13]) );
  FD_EN_55 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[14]) );
  FD_EN_54 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[15]) );
  FD_EN_53 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[16]) );
  FD_EN_52 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[17]) );
  FD_EN_51 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[18]) );
  FD_EN_50 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[19]) );
  FD_EN_49 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[20]) );
  FD_EN_48 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[21]) );
  FD_EN_47 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[22]) );
  FD_EN_46 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[23]) );
  FD_EN_45 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[24]) );
  FD_EN_44 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[25]) );
  FD_EN_43 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[26]) );
  FD_EN_42 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[27]) );
  FD_EN_41 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[28]) );
  FD_EN_40 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[29]) );
  FD_EN_39 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[30]) );
  FD_EN_38 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[31]) );
endmodule


module RegEn_Nbit32_1 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;


  FD_EN_37 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_36 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_35 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_34 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_33 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
  FD_EN_32 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[5]) );
  FD_EN_31 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[6]) );
  FD_EN_30 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[7]) );
  FD_EN_29 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[8]) );
  FD_EN_28 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[9]) );
  FD_EN_27 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[10]) );
  FD_EN_26 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[11]) );
  FD_EN_25 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[12]) );
  FD_EN_24 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[13]) );
  FD_EN_23 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[14]) );
  FD_EN_22 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[15]) );
  FD_EN_21 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[16]) );
  FD_EN_20 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[17]) );
  FD_EN_19 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[18]) );
  FD_EN_18 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[19]) );
  FD_EN_17 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[20]) );
  FD_EN_16 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[21]) );
  FD_EN_15 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[22]) );
  FD_EN_14 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[23]) );
  FD_EN_13 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[24]) );
  FD_EN_12 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[25]) );
  FD_EN_11 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[26]) );
  FD_EN_10 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[27]) );
  FD_EN_9 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[28]) );
  FD_EN_8 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[29]) );
  FD_EN_7 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[30]) );
  FD_EN_6 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[31]) );
endmodule


module FD_EN_427 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_426 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_425 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_424 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_423 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_422 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_421 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_420 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_419 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_418 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_417 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_416 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_415 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_414 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_413 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_412 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_411 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_410 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_409 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_408 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_407 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_406 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_405 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_404 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_403 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_402 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_401 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_400 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_399 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_398 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_397 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_396 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_395 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_394 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_393 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_392 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_391 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_390 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_389 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_388 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_387 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_386 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_385 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_384 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_383 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_382 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_381 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_380 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_371 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n21) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
endmodule


module FD_EN_370 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n21) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
endmodule


module FD_EN_369 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n21) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
endmodule


module FD_EN_368 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n21) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
endmodule


module FD_EN_367 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_366 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_365 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_364 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_363 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_362 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_361 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_360 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_359 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_358 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_357 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_356 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_355 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_354 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_353 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_352 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_351 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_350 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_349 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_348 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_347 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_346 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_345 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_344 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_343 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_342 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_341 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_340 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_339 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_338 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_337 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_336 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_335 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_334 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_333 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_332 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_331 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_330 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_329 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_328 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_327 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_326 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_325 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_324 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_323 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_322 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_321 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_320 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_319 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_318 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_317 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_316 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_315 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_314 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_313 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_312 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_311 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_310 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_309 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_308 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_307 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_306 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_305 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_304 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_303 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_302 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_301 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_300 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_299 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_298 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_297 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_296 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_295 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_294 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_293 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_292 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_291 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_290 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_289 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_288 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_287 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_286 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_285 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_284 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_283 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_282 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_281 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_280 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_279 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_278 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_277 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_276 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_275 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_274 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_273 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_272 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_271 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_270 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_269 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_268 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_267 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_266 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_265 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_264 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_263 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_262 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_261 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_260 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_259 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_258 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_257 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_256 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_255 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_254 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_253 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_252 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_251 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_250 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_249 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_248 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_247 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_246 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_245 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_244 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_243 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_242 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_241 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_240 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;
  tri   D;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_239 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_238 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_237 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_236 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_235 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_234 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_233 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_232 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_231 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_230 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_229 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_228 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_227 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_226 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_225 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_224 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_223 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_222 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_221 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_220 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_219 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_218 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_217 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_216 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_215 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_214 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_213 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_212 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_211 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_210 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_209 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_208 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_207 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_206 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_205 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_204 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_203 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_202 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_201 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_200 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_199 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_198 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_197 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_196 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_195 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_194 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_193 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_192 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_191 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_190 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_189 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_188 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_187 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_186 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_185 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_184 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_183 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_182 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_181 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_180 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_179 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_178 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_177 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_176 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_175 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_174 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_173 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_172 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_171 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_170 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_169 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_168 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_167 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_166 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_165 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_164 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_163 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_162 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_161 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_160 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_159 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_158 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_157 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_156 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_155 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_154 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_153 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_152 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_151 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_150 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_149 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_148 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_147 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_146 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_145 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_144 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_143 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_142 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_141 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_140 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_139 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_138 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_137 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_136 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_135 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_134 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_133 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_132 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_131 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_130 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_129 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_128 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_127 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_126 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_125 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_124 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_123 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_122 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_121 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_120 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_119 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_118 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_117 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_116 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_115 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_114 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_113 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_112 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_111 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_110 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_109 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_108 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_107 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_106 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_105 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_104 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_103 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_102 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_101 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_100 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_99 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_98 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_97 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_96 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_95 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_94 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_93 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_92 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_91 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_90 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_89 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_88 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_87 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_86 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_85 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_84 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_83 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_82 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_81 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_80 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_79 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_78 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_77 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_76 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_75 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_74 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_73 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_72 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_71 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_70 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_69 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_68 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_67 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_66 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_65 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_64 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_63 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_62 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_61 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_60 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_59 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_58 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_57 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_56 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_55 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_54 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_53 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_52 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_51 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_50 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_49 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_48 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_47 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_46 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_45 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_44 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_43 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_42 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_41 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_40 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_39 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_38 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_37 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_36 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_35 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_34 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_33 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_32 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_31 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_30 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_29 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_28 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_27 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_26 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_25 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_24 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_23 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_22 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_21 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_20 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_19 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_18 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_17 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_16 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_15 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_14 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_13 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_12 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_11 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_10 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_9 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_8 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_7 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_6 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_5 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_4 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_3 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_2 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module FD_EN_1 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n21, n22;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n22), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n21), .B2(Q), .ZN(n22) );
  INV_X1 U5 ( .A(EN), .ZN(n21) );
endmodule


module MUX21_52 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n15, n16;

  INV_X1 U1 ( .A(n16), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n16) );
  INV_X1 U3 ( .A(S), .ZN(n15) );
endmodule


module MUX21_362 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_361 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_360 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_359 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_358 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_118 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_117 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_115 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_114 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_113 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_112 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_110 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_109 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_108 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_107 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_105 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_104 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_103 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_102 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_100 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_99 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_98 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_97 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_95 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_94 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_93 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_92 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_90 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_89 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_88 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_87 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_85 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_84 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_83 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_82 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_47 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_791 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_790 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_789 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_788 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_787 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_786 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_785 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_784 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_783 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_782 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_781 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_780 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_779 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_778 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_777 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_776 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_775 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_774 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_773 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_772 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_771 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_770 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_769 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_768 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_766 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_765 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_764 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_763 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_762 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_761 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_760 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_759 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_758 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_757 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_756 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_755 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_754 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_753 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_752 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_751 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_750 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_749 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_748 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_747 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_746 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_745 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_744 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_743 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_742 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_741 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_740 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_739 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_738 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_737 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_736 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_734 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_733 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_732 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_731 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_730 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_729 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_728 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_727 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_726 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_725 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_724 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_723 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_722 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_721 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_720 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_719 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_718 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_717 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_716 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_715 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_714 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_713 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_712 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_711 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_710 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_709 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_708 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_707 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_706 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_705 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_704 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_700 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_699 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_698 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_697 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_696 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_695 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_694 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_693 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_692 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_691 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_690 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_689 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_688 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_687 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_686 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_685 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_684 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_683 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_682 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_681 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_680 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_679 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_678 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_677 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_676 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_675 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_674 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_673 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_672 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_671 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_670 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_669 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_668 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_667 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_666 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_665 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_664 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_663 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_662 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_661 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_660 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_659 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_658 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_657 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_656 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_655 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_654 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_653 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_652 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_651 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_650 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_649 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_647 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_646 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_645 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_644 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_643 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_642 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_641 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_640 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_639 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_638 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_637 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_636 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_635 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_634 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_633 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_632 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_631 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_630 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_629 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_628 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_627 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_626 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_625 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_624 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_623 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_622 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_621 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_620 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_619 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_618 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_617 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_616 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_615 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_614 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_613 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_612 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_611 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_610 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_609 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_608 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_607 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_606 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_605 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_604 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_603 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_602 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_601 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_600 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_599 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_598 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_597 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_596 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_595 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_594 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_593 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_592 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_591 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_590 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_589 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_588 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_587 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_586 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_585 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_584 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_583 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_582 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_581 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_580 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_579 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_578 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_577 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_566 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_565 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_564 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_563 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_562 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_561 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_560 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_559 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_558 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_557 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_556 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_555 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_554 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_553 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_552 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_551 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_550 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_549 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_548 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_547 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_546 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_545 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_544 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_543 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_542 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_541 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_540 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_539 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_538 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_537 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_536 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_535 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;
  tri   in1;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_534 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_533 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_532 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_531 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_530 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_529 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_528 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_527 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_526 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_525 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_524 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_523 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_522 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_521 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_520 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_519 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_518 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_517 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_516 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_515 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_514 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_513 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_512 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_511 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_510 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_509 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_508 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_507 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_506 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_505 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_504 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_503 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_500 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_496 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_492 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_490 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_489 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_488 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_487 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_485 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_484 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_483 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_482 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_481 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_480 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_478 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_477 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_476 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_475 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_474 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_473 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_472 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_471 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_470 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_468 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_467 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_466 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_465 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_464 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_463 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_462 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_461 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_460 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_459 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_458 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_457 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_456 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_455 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_454 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_453 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_452 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_451 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_450 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_449 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_448 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_447 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_446 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_445 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_444 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_443 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_442 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_441 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_440 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_439 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_431 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_430 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_429 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_428 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_427 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_426 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_425 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_424 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_423 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_422 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_421 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_420 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_419 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_418 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_417 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_416 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_415 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_414 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_413 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_412 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_411 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_410 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_409 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_408 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_407 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_406 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_405 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_404 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_403 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_402 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_401 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_400 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_399 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_398 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_397 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_396 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_395 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_394 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_393 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_392 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_391 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_390 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_389 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_388 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_387 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_386 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_385 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_384 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_383 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_382 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_381 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_380 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_379 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_378 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_377 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_376 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_375 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_374 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_373 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_372 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_371 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_370 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_369 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_368 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_326 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_325 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_321 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_295 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  AOI22_X1 U1 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U2 ( .A(S), .ZN(n16) );
  INV_X1 U3 ( .A(n17), .ZN(Y) );
endmodule


module MUX21_293 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  AOI22_X1 U1 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U2 ( .A(S), .ZN(n16) );
  INV_X1 U3 ( .A(n17), .ZN(Y) );
endmodule


module MUX21_291 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_290 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_289 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_80 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_79 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_78 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_77 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_76 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n16, n17;

  INV_X1 U1 ( .A(n17), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n17) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_571 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_570 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_569 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_568 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_567 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_495 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_357 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_356 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_355 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_354 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_353 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_265 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_263 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_262 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_261 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_260 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_259 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_258 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_257 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_256 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_255 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_254 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_253 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_252 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_251 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_250 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_249 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_248 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_247 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_246 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_245 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_244 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_243 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_242 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_241 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_240 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_239 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_238 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_237 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_236 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_235 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_234 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_233 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_232 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_231 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_230 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_229 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_228 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_227 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_226 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_225 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_224 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_223 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_222 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_221 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_220 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_219 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_218 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_217 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_216 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_215 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_214 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_213 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_212 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_211 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_210 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_209 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_208 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_207 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_206 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_205 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_204 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_203 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_202 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_201 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_200 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_199 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_198 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_197 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_196 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_195 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_194 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_193 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_192 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_191 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_190 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_189 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_188 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_187 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_186 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_185 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_184 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_183 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_182 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_181 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_180 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_179 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_178 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_177 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_176 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_175 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_174 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_173 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_172 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_171 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_170 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_169 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_168 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_167 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_166 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_165 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_164 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_163 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_162 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_161 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_160 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_159 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_158 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_157 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_156 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_152 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_151 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_146 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_141 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_136 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_131 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_126 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_121 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_120 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_119 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n18), .ZN(Y) );
endmodule


module MUX21_116 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_111 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_106 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_101 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_96 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_91 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_86 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_81 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_75 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_74 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_73 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_70 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_61 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_60 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_46 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_275 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_155 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_154 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_153 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_150 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_149 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_148 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_147 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_145 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_144 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_143 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_142 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_140 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_139 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_138 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_137 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
  INV_X1 U3 ( .A(S), .ZN(n17) );
endmodule


module MUX21_135 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_134 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_133 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_132 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_129 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_128 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_127 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_125 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_124 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_123 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_122 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  INV_X1 U2 ( .A(n18), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_71 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_66 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_56 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_51 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module MUX21_41 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n17, n18;

  INV_X1 U1 ( .A(n18), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  AOI22_X1 U3 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n18) );
endmodule


module RCAN_Nbit4_55 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_667 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_666 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_665 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_664 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_54 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_663 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_662 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_661 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_660 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_53 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_659 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_658 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_657 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_656 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_52 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_655 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_654 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_653 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_652 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_51 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_651 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_650 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_649 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_648 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_50 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_647 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_646 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_645 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_644 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_49 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_643 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_642 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_641 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_640 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_46 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_631 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_630 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_629 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_628 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_45 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_627 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_626 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_625 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_624 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_44 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_623 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_622 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_621 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_620 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_43 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_619 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_618 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_617 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_616 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_42 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_615 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_614 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_613 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_612 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_41 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_611 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_610 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_609 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_608 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_40 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_607 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_606 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_605 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_604 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_39 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_603 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_602 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_601 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_600 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_38 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_599 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_598 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_597 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_596 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_37 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_595 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_594 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_593 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_592 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_36 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_591 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_590 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_589 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_588 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_35 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_587 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_586 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_585 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_584 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_34 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_583 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_582 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_581 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_580 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_33 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_579 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_578 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_577 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_576 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_32 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_575 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_574 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_573 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_572 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_45 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n9, n10;

  AOI22_X1 U1 ( .A1(n9), .A2(in0), .B1(S), .B2(in1), .ZN(n10) );
  INV_X1 U2 ( .A(S), .ZN(n9) );
  INV_X1 U3 ( .A(n10), .ZN(Y) );
endmodule


module PG_42 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n7;

  INV_X1 U1 ( .A(n7), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n7) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module MUX21_266 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n15, n16;
  tri   S;

  INV_X1 U1 ( .A(n16), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n15) );
  AOI22_X1 U3 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n16) );
endmodule


module MUX21_67 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n15, n16;

  INV_X1 U1 ( .A(n16), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n16) );
  INV_X1 U3 ( .A(S), .ZN(n15) );
endmodule


module MUX21_62 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n15, n16;

  INV_X1 U1 ( .A(n16), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n16) );
  INV_X1 U3 ( .A(S), .ZN(n15) );
endmodule


module MUX21_53 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n15, n16;

  INV_X1 U1 ( .A(n16), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n16) );
  INV_X1 U3 ( .A(S), .ZN(n15) );
endmodule


module MUX21_267 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n15, n16;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n15) );
  INV_X1 U2 ( .A(n16), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n16) );
endmodule


module MUX21_130 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n9, n10;

  INV_X1 U1 ( .A(S), .ZN(n9) );
  INV_X1 U2 ( .A(n10), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n9), .B1(in1), .B2(S), .ZN(n10) );
endmodule


module MUX21_44 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n11, n12;

  AOI22_X1 U1 ( .A1(in0), .A2(n11), .B1(S), .B2(in1), .ZN(n12) );
  INV_X1 U2 ( .A(S), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
endmodule


module FA_560 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n18), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n18) );
  INV_X1 U1 ( .A(n17), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n18), .B2(Ci), .ZN(n17) );
endmodule


module FA_549 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n18), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n18) );
  INV_X1 U1 ( .A(n17), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n18), .B2(Ci), .ZN(n17) );
endmodule


module FA_547 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n18), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n18) );
  INV_X1 U1 ( .A(n17), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n18), .B2(Ci), .ZN(n17) );
endmodule


module FA_527 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n17, n18;

  XOR2_X1 U3 ( .A(Ci), .B(n18), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n18) );
  INV_X1 U1 ( .A(n17), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n18), .B2(Ci), .ZN(n17) );
endmodule


module MUX21_42 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n13, n14;

  AOI22_X1 U1 ( .A1(in0), .A2(n13), .B1(S), .B2(in1), .ZN(n14) );
  INV_X1 U2 ( .A(S), .ZN(n13) );
  INV_X1 U3 ( .A(n14), .ZN(Y) );
endmodule


module FD_EN_379 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n15, n16;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n15) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n16), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n15), .B2(Q), .ZN(n16) );
endmodule


module FD_EN_374 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n15, n16;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n15) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n16), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n15), .B2(Q), .ZN(n16) );
endmodule


module MUX21_469 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n10, n11;

  INV_X1 U1 ( .A(n11), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n11) );
  INV_X1 U3 ( .A(S), .ZN(n10) );
endmodule


module MUX21_433 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n10, n11;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n10) );
  INV_X1 U2 ( .A(n11), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n11) );
endmodule


module MUX21_273 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n10, n11;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n10) );
  AOI22_X1 U2 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n11) );
  INV_X1 U3 ( .A(n11), .ZN(Y) );
endmodule


module MUX21_57 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n10, n11;

  INV_X1 U1 ( .A(n11), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n11) );
  INV_X1 U3 ( .A(S), .ZN(n10) );
endmodule


module mux21N_N5_32 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_160 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_159 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_158 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_157 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_156 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module MUX21_1 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_2 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_3 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_4 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_5 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_6 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_7 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_8 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_9 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_10 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_11 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_12 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_13 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_14 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_15 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_16 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_17 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_18 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_19 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_20 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_21 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_22 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_23 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_24 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_25 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_26 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_27 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_28 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_29 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_30 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_31 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_32 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_33 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_34 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_35 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Co) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Co) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_36 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_37 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_38 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_39 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_0 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Co) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Co) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_0_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_43 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module FA_515 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_516 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_519 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_48 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_49 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(S), .B2(in1), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_50 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(S), .B2(in1), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module FA_520 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_522 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_523 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_524 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_525 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_54 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_55 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module FA_531 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_535 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_58 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_59 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module FA_536 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_537 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_538 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Co) );
endmodule


module FA_539 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_540 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_541 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_543 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_63 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_64 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_65 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module FA_544 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_546 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_551 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_68 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_69 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module FA_552 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_553 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_554 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_555 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n2) );
  CLKBUF_X1 U1 ( .A(B), .Z(n15) );
  INV_X1 U2 ( .A(n3), .ZN(Co) );
  AOI22_X1 U5 ( .A1(n15), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_556 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_558 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_559 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_72 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module FA_562 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_563 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_564 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_565 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_566 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_567 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_570 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_571 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module mux21N_N5_1 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;
  wire   n2;
  assign n2 = S;

  MUX21_5 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n2), .Y(U[0]) );
  MUX21_4 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n2), .Y(U[1]) );
  MUX21_3 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n2), .Y(U[2]) );
  MUX21_2 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n2), .Y(U[3]) );
  MUX21_1 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n2), .Y(U[4]) );
endmodule


module RCAN_Nbit4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(CTMP_2_port) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(CTMP_3_port) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(CTMP_2_port) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(CTMP_3_port) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_2 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;
  wire   n2;
  assign n2 = S;

  MUX21_10 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n2), .Y(U[0]) );
  MUX21_9 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n2), .Y(U[1]) );
  MUX21_8 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n2), .Y(U[2]) );
  MUX21_7 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n2), .Y(U[3]) );
  MUX21_6 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n2), .Y(U[4]) );
endmodule


module RCAN_Nbit4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_3 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_15 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_14 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_13 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_12 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_11 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_4 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_20 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_19 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_18 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_17 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_16 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_5 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_25 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_24 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_23 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_22 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_21 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_6 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_30 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_29 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_28 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_27 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_26 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_7 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_35 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_34 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_33 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_32 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_31 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_0 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_0 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_39 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_38 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_37 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_36 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   CTMP_1_port, CTMP_2_port, CTMP_3_port;

  FA_0_1 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP_1_port) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP_1_port), .S(S[1]), .Co(
        CTMP_2_port) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP_2_port), .S(S[2]), .Co(
        CTMP_3_port) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP_3_port), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_9 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;
  wire   n8, n9, n10;
  assign n8 = S;

  MUX21_45 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n8), .Y(U[0]) );
  MUX21_44 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n8), .Y(U[1]) );
  MUX21_43 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n8), .Y(U[2]) );
  MUX21_42 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n9), .Y(U[3]) );
  MUX21_41 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n10), .Y(U[4]) );
  BUF_X1 U1 ( .A(n8), .Z(n9) );
  CLKBUF_X1 U2 ( .A(n9), .Z(n10) );
endmodule


module RCAN_Nbit4_17 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_515 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_514 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_513 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_512 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_18 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_519 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_518 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_517 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_516 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_10 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;
  wire   n6, n7;
  assign n6 = S;

  MUX21_50 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n6), .Y(U[0]) );
  MUX21_49 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n6), .Y(U[1]) );
  MUX21_48 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n6), .Y(U[2]) );
  MUX21_47 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n6), .Y(U[3]) );
  MUX21_46 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n7), .Y(U[4]) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n7) );
endmodule


module RCAN_Nbit4_19 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_523 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_522 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_521 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_520 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_20 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_527 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_526 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_525 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_524 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_11 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;
  wire   n6;
  assign n6 = S;

  MUX21_55 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n6), .Y(U[0]) );
  MUX21_54 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n6), .Y(U[1]) );
  MUX21_53 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n6), .Y(U[2]) );
  MUX21_52 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n6), .Y(U[3]) );
  MUX21_51 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n6), .Y(U[4]) );
endmodule


module RCAN_Nbit4_21 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_531 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_530 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_529 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_528 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_22 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_535 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_534 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_533 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_532 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_12 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;
  wire   n7;
  assign n7 = S;

  MUX21_60 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n7), .Y(U[0]) );
  MUX21_59 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n7), .Y(U[1]) );
  MUX21_58 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n7), .Y(U[2]) );
  MUX21_57 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n7), .Y(U[3]) );
  MUX21_56 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n7), .Y(U[4]) );
endmodule


module RCAN_Nbit4_23 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_539 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_538 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_537 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_536 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_24 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_543 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_542 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_541 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_540 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_13 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;
  wire   n2;
  assign n2 = S;

  MUX21_65 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n2), .Y(U[0]) );
  MUX21_64 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n2), .Y(U[1]) );
  MUX21_63 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n2), .Y(U[2]) );
  MUX21_62 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n2), .Y(U[3]) );
  MUX21_61 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n2), .Y(U[4]) );
endmodule


module RCAN_Nbit4_25 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_547 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_546 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_545 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_544 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_26 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_551 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_550 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_549 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_548 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_14 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;
  wire   n2;
  assign n2 = S;

  MUX21_70 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n2), .Y(U[0]) );
  MUX21_69 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n2), .Y(U[1]) );
  MUX21_68 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n2), .Y(U[2]) );
  MUX21_67 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n2), .Y(U[3]) );
  MUX21_66 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n2), .Y(U[4]) );
endmodule


module RCAN_Nbit4_27 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_555 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_554 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_553 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_552 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_28 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_559 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_558 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_557 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_556 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_15 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_75 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_74 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_73 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_72 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_71 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_29 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_563 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_562 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_561 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_560 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_30 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_567 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_566 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_565 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_564 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_16 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_80 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_79 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_78 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_77 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_76 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_31 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_571 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_570 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_569 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_568 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSBlockNBM_Nbit4_1 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;
  wire   sum_cin0_0_port, sum_cin0_1_port, sum_cin0_2_port, sum_cin0_3_port,
         sum_cin0_4_port, sum_cin1_0_port, sum_cin1_1_port, sum_cin1_2_port,
         sum_cin1_3_port, sum_cin1_4_port;

  RCAN_Nbit4_2 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S({sum_cin0_3_port, 
        sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), .Co(
        sum_cin0_4_port) );
  RCAN_Nbit4_1 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S({sum_cin1_3_port, 
        sum_cin1_2_port, sum_cin1_1_port, sum_cin1_0_port}), .Co(
        sum_cin1_4_port) );
  mux21N_N5_1 MUX ( .in1({sum_cin1_4_port, sum_cin1_3_port, sum_cin1_2_port, 
        sum_cin1_1_port, sum_cin1_0_port}), .in0({sum_cin0_4_port, 
        sum_cin0_3_port, sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), 
        .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockNBM_Nbit4_2 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;
  wire   sum_cin0_0_port, sum_cin0_1_port, sum_cin0_2_port, sum_cin0_3_port,
         sum_cin0_4_port, sum_cin1_0_port, sum_cin1_1_port, sum_cin1_2_port,
         sum_cin1_3_port, sum_cin1_4_port;

  RCAN_Nbit4_4 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S({sum_cin0_3_port, 
        sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), .Co(
        sum_cin0_4_port) );
  RCAN_Nbit4_3 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S({sum_cin1_3_port, 
        sum_cin1_2_port, sum_cin1_1_port, sum_cin1_0_port}), .Co(
        sum_cin1_4_port) );
  mux21N_N5_2 MUX ( .in1({sum_cin1_4_port, sum_cin1_3_port, sum_cin1_2_port, 
        sum_cin1_1_port, sum_cin1_0_port}), .in0({sum_cin0_4_port, 
        sum_cin0_3_port, sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), 
        .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockNBM_Nbit4_3 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;
  wire   sum_cin0_0_port, sum_cin0_1_port, sum_cin0_2_port, sum_cin0_3_port,
         sum_cin0_4_port, sum_cin1_0_port, sum_cin1_1_port, sum_cin1_2_port,
         sum_cin1_3_port, sum_cin1_4_port;

  RCAN_Nbit4_6 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S({sum_cin0_3_port, 
        sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), .Co(
        sum_cin0_4_port) );
  RCAN_Nbit4_5 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S({sum_cin1_3_port, 
        sum_cin1_2_port, sum_cin1_1_port, sum_cin1_0_port}), .Co(
        sum_cin1_4_port) );
  mux21N_N5_3 MUX ( .in1({sum_cin1_4_port, sum_cin1_3_port, sum_cin1_2_port, 
        sum_cin1_1_port, sum_cin1_0_port}), .in0({sum_cin0_4_port, 
        sum_cin0_3_port, sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), 
        .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockNBM_Nbit4_4 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;
  wire   sum_cin0_0_port, sum_cin0_1_port, sum_cin0_2_port, sum_cin0_3_port,
         sum_cin0_4_port, sum_cin1_0_port, sum_cin1_1_port, sum_cin1_2_port,
         sum_cin1_3_port, sum_cin1_4_port;

  RCAN_Nbit4_8 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S({sum_cin0_3_port, 
        sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), .Co(
        sum_cin0_4_port) );
  RCAN_Nbit4_7 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S({sum_cin1_3_port, 
        sum_cin1_2_port, sum_cin1_1_port, sum_cin1_0_port}), .Co(
        sum_cin1_4_port) );
  mux21N_N5_4 MUX ( .in1({sum_cin1_4_port, sum_cin1_3_port, sum_cin1_2_port, 
        sum_cin1_1_port, sum_cin1_0_port}), .in0({sum_cin0_4_port, 
        sum_cin0_3_port, sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), 
        .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockNBM_Nbit4_5 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;
  wire   sum_cin0_0_port, sum_cin0_1_port, sum_cin0_2_port, sum_cin0_3_port,
         sum_cin0_4_port, sum_cin1_0_port, sum_cin1_1_port, sum_cin1_2_port,
         sum_cin1_3_port, sum_cin1_4_port;

  RCAN_Nbit4_10 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S({sum_cin0_3_port, 
        sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), .Co(
        sum_cin0_4_port) );
  RCAN_Nbit4_9 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S({sum_cin1_3_port, 
        sum_cin1_2_port, sum_cin1_1_port, sum_cin1_0_port}), .Co(
        sum_cin1_4_port) );
  mux21N_N5_5 MUX ( .in1({sum_cin1_4_port, sum_cin1_3_port, sum_cin1_2_port, 
        sum_cin1_1_port, sum_cin1_0_port}), .in0({sum_cin0_4_port, 
        sum_cin0_3_port, sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), 
        .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockNBM_Nbit4_6 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;
  wire   sum_cin0_0_port, sum_cin0_1_port, sum_cin0_2_port, sum_cin0_3_port,
         sum_cin0_4_port, sum_cin1_0_port, sum_cin1_1_port, sum_cin1_2_port,
         sum_cin1_3_port, sum_cin1_4_port;

  RCAN_Nbit4_12 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S({sum_cin0_3_port, 
        sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), .Co(
        sum_cin0_4_port) );
  RCAN_Nbit4_11 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S({sum_cin1_3_port, 
        sum_cin1_2_port, sum_cin1_1_port, sum_cin1_0_port}), .Co(
        sum_cin1_4_port) );
  mux21N_N5_6 MUX ( .in1({sum_cin1_4_port, sum_cin1_3_port, sum_cin1_2_port, 
        sum_cin1_1_port, sum_cin1_0_port}), .in0({sum_cin0_4_port, 
        sum_cin0_3_port, sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), 
        .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockNBM_Nbit4_7 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;
  wire   sum_cin0_0_port, sum_cin0_1_port, sum_cin0_2_port, sum_cin0_3_port,
         sum_cin0_4_port, sum_cin1_0_port, sum_cin1_1_port, sum_cin1_2_port,
         sum_cin1_3_port, sum_cin1_4_port;

  RCAN_Nbit4_14 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S({sum_cin0_3_port, 
        sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), .Co(
        sum_cin0_4_port) );
  RCAN_Nbit4_13 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S({sum_cin1_3_port, 
        sum_cin1_2_port, sum_cin1_1_port, sum_cin1_0_port}), .Co(
        sum_cin1_4_port) );
  mux21N_N5_7 MUX ( .in1({sum_cin1_4_port, sum_cin1_3_port, sum_cin1_2_port, 
        sum_cin1_1_port, sum_cin1_0_port}), .in0({sum_cin0_4_port, 
        sum_cin0_3_port, sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), 
        .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockNBM_Nbit4_0 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;
  wire   sum_cin0_0_port, sum_cin0_1_port, sum_cin0_2_port, sum_cin0_3_port,
         sum_cin0_4_port, sum_cin1_0_port, sum_cin1_1_port, sum_cin1_2_port,
         sum_cin1_3_port, sum_cin1_4_port;

  RCAN_Nbit4_0 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S({sum_cin0_3_port, 
        sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), .Co(
        sum_cin0_4_port) );
  RCAN_Nbit4_15 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S({sum_cin1_3_port, 
        sum_cin1_2_port, sum_cin1_1_port, sum_cin1_0_port}), .Co(
        sum_cin1_4_port) );
  mux21N_N5_0 MUX ( .in1({sum_cin1_4_port, sum_cin1_3_port, sum_cin1_2_port, 
        sum_cin1_1_port, sum_cin1_0_port}), .in0({sum_cin0_4_port, 
        sum_cin0_3_port, sum_cin0_2_port, sum_cin0_1_port, sum_cin0_0_port}), 
        .S(Ci), .U({Cout, S}) );
endmodule


module G_1 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_2 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_3 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_4 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PG_1 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_2 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AOI21_X1 U1 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module G_5 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_6 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PG_3 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_4 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_5 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module G_7 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PG_6 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_7 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_8 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_9 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_10 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_11 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_12 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AOI21_X1 U1 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module G_8 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PG_13 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_14 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_15 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_16 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_17 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_18 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_19 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AOI21_X1 U1 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module PG_20 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_21 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_22 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_23 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_24 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_25 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_26 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_0 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AOI21_X1 U1 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module G_0 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PGblock_1 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_2 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_3 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_4 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_5 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_6 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_7 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_8 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_9 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_10 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_11 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_12 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_13 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_14 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_15 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_16 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_17 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_18 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_19 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_20 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_21 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_22 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_23 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_24 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_25 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_26 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_27 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_28 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_29 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_30 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_31 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_0 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module FA_632 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Co) );
endmodule


module FA_636 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Co) );
endmodule


module FA_694 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_695 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_696 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Co) );
endmodule


module FA_697 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_698 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_699 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_700 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Co) );
endmodule


module FA_701 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_702 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module CSBlockN_Nbit4_1 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_18 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_17 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_9 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_2 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_20 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_19 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_10 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_3 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_22 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_21 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_11 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_4 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_24 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_23 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_12 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_5 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_26 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_25 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_13 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_6 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_28 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_27 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_14 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_7 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_30 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_29 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_15 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_8 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_32 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_31 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_16 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module G_11 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   net299432, n2;
  assign Gout = net299432;

  INV_X1 U1 ( .A(n2), .ZN(net299432) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module G_12 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_13 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_29 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module G_14 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module G_15 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PG_31 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module PG_32 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module G_16 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   net396859, n2;
  assign Gout = net396859;

  INV_X1 U1 ( .A(n2), .ZN(net396859) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_33 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_34 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AOI21_X1 U1 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module PG_35 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_36 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module PG_37 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module PG_38 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_39 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module G_17 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_43 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_44 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module PG_45 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module PG_46 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PG_47 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AOI21_X1 U1 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module PG_48 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_49 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_50 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PG_51 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_52 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_53 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module PG_54 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AOI21_X1 U1 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
  AND2_X1 U2 ( .A1(P1), .A2(P2), .ZN(Pout) );
  INV_X1 U3 ( .A(n2), .ZN(Gout) );
endmodule


module G_18 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   net352122, n2;
  assign Gout = net352122;

  AOI21_X1 U1 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(net352122) );
endmodule


module PGblock_49 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_51 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_53 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_55 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_56 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_57 ( A, B, G, P );
  input A, B;
  output G, P;
  wire   n3;

  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  AND2_X1 U3 ( .A1(n3), .A2(A), .ZN(G) );
endmodule


module PGblock_61 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_63 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_64 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module CarrySumNBM_Nbit32 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  CSBlockNBM_Nbit4_0 CSN_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  CSBlockNBM_Nbit4_7 CSN_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  CSBlockNBM_Nbit4_6 CSN_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8])
         );
  CSBlockNBM_Nbit4_5 CSN_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  CSBlockNBM_Nbit4_4 CSN_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  CSBlockNBM_Nbit4_3 CSN_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  CSBlockNBM_Nbit4_2 CSN_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  CSBlockNBM_Nbit4_1 CSN_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module SparseTreeCarryGenNBM_Nbit32 ( A, B, Cin, Cout );
  input [31:0] A;
  input [31:0] B;
  output [8:0] Cout;
  input Cin;
  wire   Cin, gen_0_1_port, gen_0_2_port, prop_0_2_port, gen_0_3_port,
         prop_0_3_port, gen_0_4_port, prop_0_4_port, gen_0_5_port,
         prop_0_5_port, gen_0_6_port, prop_0_6_port, gen_0_7_port,
         prop_0_7_port, gen_0_8_port, prop_0_8_port, gen_0_9_port,
         prop_0_9_port, gen_0_10_port, prop_0_10_port, gen_0_11_port,
         prop_0_11_port, gen_0_12_port, prop_0_12_port, gen_0_13_port,
         prop_0_13_port, gen_0_14_port, prop_0_14_port, gen_0_15_port,
         prop_0_15_port, gen_0_16_port, prop_0_16_port, gen_0_17_port,
         prop_0_17_port, gen_0_18_port, prop_0_18_port, gen_0_19_port,
         prop_0_19_port, gen_0_20_port, prop_0_20_port, gen_0_21_port,
         prop_0_21_port, gen_0_22_port, prop_0_22_port, gen_0_23_port,
         prop_0_23_port, gen_0_24_port, prop_0_24_port, gen_0_25_port,
         prop_0_25_port, gen_0_26_port, prop_0_26_port, gen_0_27_port,
         prop_0_27_port, gen_0_28_port, prop_0_28_port, gen_0_29_port,
         prop_0_29_port, gen_0_30_port, prop_0_30_port, gen_0_31_port,
         prop_0_31_port, gen_0_32_port, prop_0_32_port, gen_1_2_port,
         gen_1_4_port, prop_1_4_port, gen_1_6_port, prop_1_6_port,
         gen_1_8_port, prop_1_8_port, gen_1_10_port, prop_1_10_port,
         gen_1_12_port, prop_1_12_port, gen_1_14_port, prop_1_14_port,
         gen_1_16_port, prop_1_16_port, gen_1_18_port, prop_1_18_port,
         gen_1_20_port, prop_1_20_port, gen_1_22_port, prop_1_22_port,
         gen_1_24_port, prop_1_24_port, gen_1_26_port, prop_1_26_port,
         gen_1_28_port, prop_1_28_port, gen_1_30_port, prop_1_30_port,
         gen_1_32_port, prop_1_32_port, gen_2_8_port, prop_2_8_port,
         gen_2_12_port, prop_2_12_port, gen_2_16_port, prop_2_16_port,
         prop_2_20_port, gen_2_24_port, prop_2_24_port, gen_2_28_port,
         prop_2_28_port, gen_2_32_port, prop_2_32_port, gen_3_16_port,
         prop_3_16_port, prop_3_24_port, gen_3_32_port, prop_3_32_port,
         gen_4_28_port, prop_4_28_port, n3, gen_4_32_port, prop_4_32_port, n2;
  assign Cout[0] = Cin;

  PGblock_0 PGB_0_1 ( .A(A[0]), .B(B[0]), .G(gen_0_1_port) );
  PGblock_31 PGB_0_2 ( .A(A[1]), .B(B[1]), .G(gen_0_2_port), .P(prop_0_2_port)
         );
  PGblock_30 PGB_0_3 ( .A(A[2]), .B(B[2]), .G(gen_0_3_port), .P(prop_0_3_port)
         );
  PGblock_29 PGB_0_4 ( .A(A[3]), .B(B[3]), .G(gen_0_4_port), .P(prop_0_4_port)
         );
  PGblock_28 PGB_0_5 ( .A(A[4]), .B(B[4]), .G(gen_0_5_port), .P(prop_0_5_port)
         );
  PGblock_27 PGB_0_6 ( .A(A[5]), .B(B[5]), .G(gen_0_6_port), .P(prop_0_6_port)
         );
  PGblock_26 PGB_0_7 ( .A(A[6]), .B(B[6]), .G(gen_0_7_port), .P(prop_0_7_port)
         );
  PGblock_25 PGB_0_8 ( .A(A[7]), .B(B[7]), .G(gen_0_8_port), .P(prop_0_8_port)
         );
  PGblock_24 PGB_0_9 ( .A(A[8]), .B(B[8]), .G(gen_0_9_port), .P(prop_0_9_port)
         );
  PGblock_23 PGB_0_10 ( .A(A[9]), .B(B[9]), .G(gen_0_10_port), .P(
        prop_0_10_port) );
  PGblock_22 PGB_0_11 ( .A(A[10]), .B(B[10]), .G(gen_0_11_port), .P(
        prop_0_11_port) );
  PGblock_21 PGB_0_12 ( .A(A[11]), .B(B[11]), .G(gen_0_12_port), .P(
        prop_0_12_port) );
  PGblock_20 PGB_0_13 ( .A(A[12]), .B(B[12]), .G(gen_0_13_port), .P(
        prop_0_13_port) );
  PGblock_19 PGB_0_14 ( .A(A[13]), .B(B[13]), .G(gen_0_14_port), .P(
        prop_0_14_port) );
  PGblock_18 PGB_0_15 ( .A(A[14]), .B(B[14]), .G(gen_0_15_port), .P(
        prop_0_15_port) );
  PGblock_17 PGB_0_16 ( .A(A[15]), .B(B[15]), .G(gen_0_16_port), .P(
        prop_0_16_port) );
  PGblock_16 PGB_0_17 ( .A(A[16]), .B(B[16]), .G(gen_0_17_port), .P(
        prop_0_17_port) );
  PGblock_15 PGB_0_18 ( .A(A[17]), .B(B[17]), .G(gen_0_18_port), .P(
        prop_0_18_port) );
  PGblock_14 PGB_0_19 ( .A(A[18]), .B(B[18]), .G(gen_0_19_port), .P(
        prop_0_19_port) );
  PGblock_13 PGB_0_20 ( .A(A[19]), .B(B[19]), .G(gen_0_20_port), .P(
        prop_0_20_port) );
  PGblock_12 PGB_0_21 ( .A(A[20]), .B(B[20]), .G(gen_0_21_port), .P(
        prop_0_21_port) );
  PGblock_11 PGB_0_22 ( .A(A[21]), .B(B[21]), .G(gen_0_22_port), .P(
        prop_0_22_port) );
  PGblock_10 PGB_0_23 ( .A(A[22]), .B(B[22]), .G(gen_0_23_port), .P(
        prop_0_23_port) );
  PGblock_9 PGB_0_24 ( .A(A[23]), .B(B[23]), .G(gen_0_24_port), .P(
        prop_0_24_port) );
  PGblock_8 PGB_0_25 ( .A(A[24]), .B(B[24]), .G(gen_0_25_port), .P(
        prop_0_25_port) );
  PGblock_7 PGB_0_26 ( .A(A[25]), .B(B[25]), .G(gen_0_26_port), .P(
        prop_0_26_port) );
  PGblock_6 PGB_0_27 ( .A(A[26]), .B(B[26]), .G(gen_0_27_port), .P(
        prop_0_27_port) );
  PGblock_5 PGB_0_28 ( .A(A[27]), .B(B[27]), .G(gen_0_28_port), .P(
        prop_0_28_port) );
  PGblock_4 PGB_0_29 ( .A(A[28]), .B(B[28]), .G(gen_0_29_port), .P(
        prop_0_29_port) );
  PGblock_3 PGB_0_30 ( .A(A[29]), .B(B[29]), .G(gen_0_30_port), .P(
        prop_0_30_port) );
  PGblock_2 PGB_0_31 ( .A(A[30]), .B(B[30]), .G(gen_0_31_port), .P(
        prop_0_31_port) );
  PGblock_1 PGB_0_32 ( .A(A[31]), .B(B[31]), .G(gen_0_32_port), .P(
        prop_0_32_port) );
  G_0 G1_2_1_1 ( .G1(gen_0_2_port), .P1(prop_0_2_port), .G2(gen_0_1_port), 
        .Gout(gen_1_2_port) );
  PG_0 PG1_2_1_2 ( .G1(gen_0_4_port), .P1(prop_0_4_port), .G2(gen_0_3_port), 
        .P2(prop_0_3_port), .Gout(gen_1_4_port), .Pout(prop_1_4_port) );
  PG_26 PG1_2_1_3 ( .G1(gen_0_6_port), .P1(prop_0_6_port), .G2(gen_0_5_port), 
        .P2(prop_0_5_port), .Gout(gen_1_6_port), .Pout(prop_1_6_port) );
  PG_25 PG1_2_1_4 ( .G1(gen_0_8_port), .P1(prop_0_8_port), .G2(gen_0_7_port), 
        .P2(prop_0_7_port), .Gout(gen_1_8_port), .Pout(prop_1_8_port) );
  PG_24 PG1_2_1_5 ( .G1(gen_0_10_port), .P1(prop_0_10_port), .G2(gen_0_9_port), 
        .P2(prop_0_9_port), .Gout(gen_1_10_port), .Pout(prop_1_10_port) );
  PG_23 PG1_2_1_6 ( .G1(gen_0_12_port), .P1(prop_0_12_port), .G2(gen_0_11_port), .P2(prop_0_11_port), .Gout(gen_1_12_port), .Pout(prop_1_12_port) );
  PG_22 PG1_2_1_7 ( .G1(gen_0_14_port), .P1(prop_0_14_port), .G2(gen_0_13_port), .P2(prop_0_13_port), .Gout(gen_1_14_port), .Pout(prop_1_14_port) );
  PG_21 PG1_2_1_8 ( .G1(gen_0_16_port), .P1(prop_0_16_port), .G2(gen_0_15_port), .P2(prop_0_15_port), .Gout(gen_1_16_port), .Pout(prop_1_16_port) );
  PG_20 PG1_2_1_9 ( .G1(gen_0_18_port), .P1(prop_0_18_port), .G2(gen_0_17_port), .P2(prop_0_17_port), .Gout(gen_1_18_port), .Pout(prop_1_18_port) );
  PG_19 PG1_2_1_10 ( .G1(gen_0_20_port), .P1(prop_0_20_port), .G2(
        gen_0_19_port), .P2(prop_0_19_port), .Gout(gen_1_20_port), .Pout(
        prop_1_20_port) );
  PG_18 PG1_2_1_11 ( .G1(gen_0_22_port), .P1(prop_0_22_port), .G2(
        gen_0_21_port), .P2(prop_0_21_port), .Gout(gen_1_22_port), .Pout(
        prop_1_22_port) );
  PG_17 PG1_2_1_12 ( .G1(gen_0_24_port), .P1(prop_0_24_port), .G2(
        gen_0_23_port), .P2(prop_0_23_port), .Gout(gen_1_24_port), .Pout(
        prop_1_24_port) );
  PG_16 PG1_2_1_13 ( .G1(gen_0_26_port), .P1(prop_0_26_port), .G2(
        gen_0_25_port), .P2(prop_0_25_port), .Gout(gen_1_26_port), .Pout(
        prop_1_26_port) );
  PG_15 PG1_2_1_14 ( .G1(gen_0_28_port), .P1(prop_0_28_port), .G2(
        gen_0_27_port), .P2(prop_0_27_port), .Gout(gen_1_28_port), .Pout(
        prop_1_28_port) );
  PG_14 PG1_2_1_15 ( .G1(gen_0_30_port), .P1(prop_0_30_port), .G2(
        gen_0_29_port), .P2(prop_0_29_port), .Gout(gen_1_30_port), .Pout(
        prop_1_30_port) );
  PG_13 PG1_2_1_16 ( .G1(gen_0_32_port), .P1(prop_0_32_port), .G2(
        gen_0_31_port), .P2(prop_0_31_port), .Gout(gen_1_32_port), .Pout(
        prop_1_32_port) );
  G_8 G1_2_2_1 ( .G1(gen_1_4_port), .P1(prop_1_4_port), .G2(gen_1_2_port), 
        .Gout(Cout[1]) );
  PG_12 PG1_2_2_2 ( .G1(gen_1_8_port), .P1(prop_1_8_port), .G2(gen_1_6_port), 
        .P2(prop_1_6_port), .Gout(gen_2_8_port), .Pout(prop_2_8_port) );
  PG_11 PG1_2_2_3 ( .G1(gen_1_12_port), .P1(prop_1_12_port), .G2(gen_1_10_port), .P2(prop_1_10_port), .Gout(gen_2_12_port), .Pout(prop_2_12_port) );
  PG_10 PG1_2_2_4 ( .G1(gen_1_16_port), .P1(prop_1_16_port), .G2(gen_1_14_port), .P2(prop_1_14_port), .Gout(gen_2_16_port), .Pout(prop_2_16_port) );
  PG_9 PG1_2_2_5 ( .G1(gen_1_20_port), .P1(prop_1_20_port), .G2(gen_1_18_port), 
        .P2(prop_1_18_port), .Gout(n2), .Pout(prop_2_20_port) );
  PG_8 PG1_2_2_6 ( .G1(gen_1_24_port), .P1(prop_1_24_port), .G2(gen_1_22_port), 
        .P2(prop_1_22_port), .Gout(gen_2_24_port), .Pout(prop_2_24_port) );
  PG_7 PG1_2_2_7 ( .G1(gen_1_28_port), .P1(prop_1_28_port), .G2(gen_1_26_port), 
        .P2(prop_1_26_port), .Gout(gen_2_28_port), .Pout(prop_2_28_port) );
  PG_6 PG1_2_2_8 ( .G1(gen_1_32_port), .P1(prop_1_32_port), .G2(gen_1_30_port), 
        .P2(prop_1_30_port), .Gout(gen_2_32_port), .Pout(prop_2_32_port) );
  G_7 G3_3_2 ( .G1(gen_2_8_port), .P1(prop_2_8_port), .G2(Cout[1]), .Gout(
        Cout[2]) );
  PG_5 PG3_3_4 ( .G1(gen_2_16_port), .P1(prop_2_16_port), .G2(gen_2_12_port), 
        .P2(prop_2_12_port), .Gout(gen_3_16_port), .Pout(prop_3_16_port) );
  PG_4 PG3_3_6 ( .G1(gen_2_24_port), .P1(prop_2_24_port), .G2(n2), .P2(
        prop_2_20_port), .Gout(n3), .Pout(prop_3_24_port) );
  PG_3 PG3_3_8 ( .G1(gen_2_32_port), .P1(prop_2_32_port), .G2(gen_2_28_port), 
        .P2(prop_2_28_port), .Gout(gen_3_32_port), .Pout(prop_3_32_port) );
  G_6 G3_E_4_2 ( .G1(gen_2_12_port), .P1(prop_2_12_port), .G2(Cout[2]), .Gout(
        Cout[3]) );
  G_5 G3_E_4_3 ( .G1(gen_3_16_port), .P1(prop_3_16_port), .G2(Cout[2]), .Gout(
        Cout[4]) );
  PG_2 PG3_E_4_6 ( .G1(gen_2_28_port), .P1(prop_2_28_port), .G2(n3), .P2(
        prop_3_24_port), .Gout(gen_4_28_port), .Pout(prop_4_28_port) );
  PG_1 PG3_E_4_7 ( .G1(gen_3_32_port), .P1(prop_3_32_port), .G2(n3), .P2(
        prop_3_24_port), .Gout(gen_4_32_port), .Pout(prop_4_32_port) );
  G_4 G3_E_5_4 ( .G1(n2), .P1(prop_2_20_port), .G2(Cout[4]), .Gout(Cout[5]) );
  G_3 G3_E_5_5 ( .G1(n3), .P1(prop_3_24_port), .G2(Cout[4]), .Gout(Cout[6]) );
  G_2 G3_E_5_6 ( .G1(gen_4_28_port), .P1(prop_4_28_port), .G2(Cout[4]), .Gout(
        Cout[7]) );
  G_1 G3_E_5_7 ( .G1(gen_4_32_port), .P1(prop_4_32_port), .G2(Cout[4]), .Gout(
        Cout[8]) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_121 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_122 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_123 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_129 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_130 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_131 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_132 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_137 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_138 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_139 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_140 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_145 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_146 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_147 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_148 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_153 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_154 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_155 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_156 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_157 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_158 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_159 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_160 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_161 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_162 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_163 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_164 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_165 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_166 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_167 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_168 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_169 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_170 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_171 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_172 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_173 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_174 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_175 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_176 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_177 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_178 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_179 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_180 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_181 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_182 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_183 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_184 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_185 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_186 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_187 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_188 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_189 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_190 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_191 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_192 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_193 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_194 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_195 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_196 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_200 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_201 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_202 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_203 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_204 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_205 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_206 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_207 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_208 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_209 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_210 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_211 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_212 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_213 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_214 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_215 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_216 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_217 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_218 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_219 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_220 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_225 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_226 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_227 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_228 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_233 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_234 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_235 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_236 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_241 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_242 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_243 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_244 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_249 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_250 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_251 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_252 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_256 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_257 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_258 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_259 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_260 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_261 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_262 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_263 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_264 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_265 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_266 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_267 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_268 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_269 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_270 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_271 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_272 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_273 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_274 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_275 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_276 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_277 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_278 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_279 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_280 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_281 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_282 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_283 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_284 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_285 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_286 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_287 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_288 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_289 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_290 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_291 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_292 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_293 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_294 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_295 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_296 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_297 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_298 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_299 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_300 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_301 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_302 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_303 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_304 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_305 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_306 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_307 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_308 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_309 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_310 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_311 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_312 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_313 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_314 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_315 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_316 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_317 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_318 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_319 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_320 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_321 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_322 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_323 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_324 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_325 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_326 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_327 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_328 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_329 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_330 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_331 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_332 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_333 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_334 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_335 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_336 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_337 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_338 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_339 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_340 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_341 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_342 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_343 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_344 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_345 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_346 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_347 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_348 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_349 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_350 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_351 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_352 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_353 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_354 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_355 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_356 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_357 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_358 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_359 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_360 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_361 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_362 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_363 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_364 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_365 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_366 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_367 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_368 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_369 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_370 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_371 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_372 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_373 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_374 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_375 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_376 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_377 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_378 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_379 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_380 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_381 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_382 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_383 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_384 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_385 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_386 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_387 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_388 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_389 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_390 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_391 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_392 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_393 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_394 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_395 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_396 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_397 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_398 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_399 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_400 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_401 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_402 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_403 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_404 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_405 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_406 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_407 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_408 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_409 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_410 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_411 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_412 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_413 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_414 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_415 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_416 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_417 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_418 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_419 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_420 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_421 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_422 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_423 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_424 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_425 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_426 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_427 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_428 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_429 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_430 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_431 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_432 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_433 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_434 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_435 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_436 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_437 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_438 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_439 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_440 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_441 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_442 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_443 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_444 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_445 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_446 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_447 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_448 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_449 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_450 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_451 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_452 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_453 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_454 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_455 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_456 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_457 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_458 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_459 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_460 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_461 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_462 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_463 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_464 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_465 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_466 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_467 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_468 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_469 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_470 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_471 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_472 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_473 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_474 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_475 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_476 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_477 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_478 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_479 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_480 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_481 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_482 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_483 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_484 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_485 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_486 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_487 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_488 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_489 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_490 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_491 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_492 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_493 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_494 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_495 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_496 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_497 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_498 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_499 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_500 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_501 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_502 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_503 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_504 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_505 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_506 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_507 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_508 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_509 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_510 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_511 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_0_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module mux21N_N5_17 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_85 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_84 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_83 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_82 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_81 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_18 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_90 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_89 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_88 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_87 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_86 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_19 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_95 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_94 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_93 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_92 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_91 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_20 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_100 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_99 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_98 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_97 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_96 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_21 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_105 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_104 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_103 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_102 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_101 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_22 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_110 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_109 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_108 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_107 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_106 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_23 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_115 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_114 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_113 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_112 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_111 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_24 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_120 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_119 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_118 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_117 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_116 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_47 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_635 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_634 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_633 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_632 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_48 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_639 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_638 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_637 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_636 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_25 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_125 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_124 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_123 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_122 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_121 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_26 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_130 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_129 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_128 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_127 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_126 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_27 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_135 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_134 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_133 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_132 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_131 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_28 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_140 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_139 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_138 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_137 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_136 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_56 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_671 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_670 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_669 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_668 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_29 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_145 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_144 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_143 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_142 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_141 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_57 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_675 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_674 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_673 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_672 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_58 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_679 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_678 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_677 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_676 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_30 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_150 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_149 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_148 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_147 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_146 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_59 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_683 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_682 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_681 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_680 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_60 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_687 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_686 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_685 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_684 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21N_N5_31 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;


  MUX21_155 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_154 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_153 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_152 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_151 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module RCAN_Nbit4_61 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_691 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_690 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_689 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_688 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_62 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_695 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_694 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_693 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_692 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_63 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_699 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_698 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_697 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_696 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCAN_Nbit4_16 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_64 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_702 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_701 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_700 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CarrySumN_Nbit32_1 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  CSBlockN_Nbit4_8 CSN_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  CSBlockN_Nbit4_7 CSN_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  CSBlockN_Nbit4_6 CSN_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8])
         );
  CSBlockN_Nbit4_5 CSN_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(S[15:12]) );
  CSBlockN_Nbit4_4 CSN_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(S[19:16]) );
  CSBlockN_Nbit4_3 CSN_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(S[23:20]) );
  CSBlockN_Nbit4_2 CSN_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(S[27:24]) );
  CSBlockN_Nbit4_1 CSN_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(S[31:28]) );
endmodule


module SparseTreeCarryGenN_Nbit32_1 ( A, B, Cin, Cout );
  input [31:0] A;
  input [31:0] B;
  output [8:0] Cout;
  input Cin;
  wire   Cin, propcin, gencin, \gen[4][28] , \gen[4][32] , \gen[3][16] ,
         \gen[3][32] , \gen[2][8] , \gen[2][16] , \gen[2][24] , \gen[2][32] ,
         \gen[1][2] , \gen[1][4] , \gen[1][6] , \gen[1][8] , \gen[1][10] ,
         \gen[1][12] , \gen[1][14] , \gen[1][16] , \gen[1][18] , \gen[1][20] ,
         \gen[1][22] , \gen[1][24] , \gen[1][26] , \gen[1][28] , \gen[1][30] ,
         \gen[1][32] , \gen[0][1] , \gen[0][2] , \gen[0][3] , \gen[0][4] ,
         \gen[0][5] , \gen[0][6] , \gen[0][7] , \gen[0][8] , \gen[0][9] ,
         \gen[0][10] , \gen[0][11] , \gen[0][12] , \gen[0][13] , \gen[0][14] ,
         \gen[0][15] , \gen[0][16] , \gen[0][17] , \gen[0][18] , \gen[0][19] ,
         \gen[0][20] , \gen[0][21] , \gen[0][22] , \gen[0][23] , \gen[0][24] ,
         \gen[0][25] , \gen[0][26] , \gen[0][27] , \gen[0][28] , \gen[0][29] ,
         \gen[0][30] , \gen[0][31] , \gen[0][32] , \prop[4][28] ,
         \prop[4][32] , \prop[3][16] , \prop[3][24] , \prop[3][32] ,
         \prop[2][8] , \prop[2][12] , \prop[2][16] , \prop[2][20] ,
         \prop[2][24] , \prop[2][28] , \prop[2][32] , \prop[1][4] ,
         \prop[1][6] , \prop[1][8] , \prop[1][10] , \prop[1][12] ,
         \prop[1][14] , \prop[1][16] , \prop[1][18] , \prop[1][20] ,
         \prop[1][22] , \prop[1][24] , \prop[1][26] , \prop[1][28] ,
         \prop[1][30] , \prop[1][32] , \prop[0][2] , \prop[0][3] ,
         \prop[0][4] , \prop[0][5] , \prop[0][6] , \prop[0][7] , \prop[0][8] ,
         \prop[0][9] , \prop[0][10] , \prop[0][11] , \prop[0][12] ,
         \prop[0][13] , \prop[0][14] , \prop[0][15] , \prop[0][16] ,
         \prop[0][17] , \prop[0][18] , \prop[0][19] , \prop[0][20] ,
         \prop[0][21] , \prop[0][22] , \prop[0][23] , \prop[0][24] ,
         \prop[0][25] , \prop[0][26] , \prop[0][27] , \prop[0][28] ,
         \prop[0][29] , \prop[0][30] , \prop[0][31] , \prop[0][32] , n74, n75,
         n78, n79, n91, n81, n92, n2, n86, n87, n89;
  assign Cout[0] = Cin;

  PGblock_64 Cinprop_0_1 ( .A(A[0]), .B(B[0]), .G(gencin), .P(propcin) );
  PGblock_63 PGB_0_2 ( .A(A[1]), .B(B[1]), .G(\gen[0][2] ), .P(\prop[0][2] )
         );
  PGblock_62 PGB_0_3 ( .A(A[2]), .B(B[2]), .G(\gen[0][3] ), .P(\prop[0][3] )
         );
  PGblock_61 PGB_0_4 ( .A(A[3]), .B(B[3]), .G(\gen[0][4] ), .P(\prop[0][4] )
         );
  PGblock_60 PGB_0_5 ( .A(A[4]), .B(B[4]), .G(\gen[0][5] ), .P(\prop[0][5] )
         );
  PGblock_59 PGB_0_6 ( .A(A[5]), .B(B[5]), .G(\gen[0][6] ), .P(\prop[0][6] )
         );
  PGblock_58 PGB_0_7 ( .A(A[6]), .B(B[6]), .G(\gen[0][7] ), .P(\prop[0][7] )
         );
  PGblock_57 PGB_0_8 ( .A(A[7]), .B(B[7]), .G(\gen[0][8] ), .P(\prop[0][8] )
         );
  PGblock_56 PGB_0_9 ( .A(A[8]), .B(B[8]), .G(\gen[0][9] ), .P(\prop[0][9] )
         );
  PGblock_55 PGB_0_10 ( .A(A[9]), .B(B[9]), .G(\gen[0][10] ), .P(\prop[0][10] ) );
  PGblock_54 PGB_0_11 ( .A(A[10]), .B(B[10]), .G(\gen[0][11] ), .P(
        \prop[0][11] ) );
  PGblock_53 PGB_0_12 ( .A(A[11]), .B(B[11]), .G(\gen[0][12] ), .P(
        \prop[0][12] ) );
  PGblock_52 PGB_0_13 ( .A(A[12]), .B(B[12]), .G(\gen[0][13] ), .P(
        \prop[0][13] ) );
  PGblock_51 PGB_0_14 ( .A(A[13]), .B(B[13]), .G(\gen[0][14] ), .P(
        \prop[0][14] ) );
  PGblock_50 PGB_0_15 ( .A(A[14]), .B(B[14]), .G(\gen[0][15] ), .P(
        \prop[0][15] ) );
  PGblock_49 PGB_0_16 ( .A(A[15]), .B(B[15]), .G(\gen[0][16] ), .P(
        \prop[0][16] ) );
  PGblock_48 PGB_0_17 ( .A(A[16]), .B(B[16]), .G(\gen[0][17] ), .P(
        \prop[0][17] ) );
  PGblock_47 PGB_0_18 ( .A(A[17]), .B(B[17]), .G(\gen[0][18] ), .P(
        \prop[0][18] ) );
  PGblock_46 PGB_0_19 ( .A(A[18]), .B(B[18]), .G(\gen[0][19] ), .P(
        \prop[0][19] ) );
  PGblock_45 PGB_0_20 ( .A(A[19]), .B(B[19]), .G(\gen[0][20] ), .P(
        \prop[0][20] ) );
  PGblock_44 PGB_0_21 ( .A(A[20]), .B(B[20]), .G(\gen[0][21] ), .P(
        \prop[0][21] ) );
  PGblock_43 PGB_0_22 ( .A(A[21]), .B(B[21]), .G(\gen[0][22] ), .P(
        \prop[0][22] ) );
  PGblock_42 PGB_0_23 ( .A(A[22]), .B(B[22]), .G(\gen[0][23] ), .P(
        \prop[0][23] ) );
  PGblock_41 PGB_0_24 ( .A(A[23]), .B(B[23]), .G(\gen[0][24] ), .P(
        \prop[0][24] ) );
  PGblock_40 PGB_0_25 ( .A(A[24]), .B(B[24]), .G(\gen[0][25] ), .P(
        \prop[0][25] ) );
  PGblock_39 PGB_0_26 ( .A(A[25]), .B(B[25]), .G(\gen[0][26] ), .P(
        \prop[0][26] ) );
  PGblock_38 PGB_0_27 ( .A(A[26]), .B(B[26]), .G(\gen[0][27] ), .P(
        \prop[0][27] ) );
  PGblock_37 PGB_0_28 ( .A(A[27]), .B(B[27]), .G(\gen[0][28] ), .P(
        \prop[0][28] ) );
  PGblock_36 PGB_0_29 ( .A(A[28]), .B(B[28]), .G(\gen[0][29] ), .P(
        \prop[0][29] ) );
  PGblock_35 PGB_0_30 ( .A(A[29]), .B(B[29]), .G(\gen[0][30] ), .P(
        \prop[0][30] ) );
  PGblock_34 PGB_0_31 ( .A(A[30]), .B(B[30]), .G(\gen[0][31] ), .P(
        \prop[0][31] ) );
  PGblock_33 PGB_0_32 ( .A(A[31]), .B(B[31]), .G(\gen[0][32] ), .P(
        \prop[0][32] ) );
  G_18 G1_2_1_1 ( .G1(\gen[0][2] ), .P1(\prop[0][2] ), .G2(\gen[0][1] ), 
        .Gout(\gen[1][2] ) );
  PG_54 PG1_2_1_2 ( .G1(\gen[0][4] ), .P1(\prop[0][4] ), .G2(\gen[0][3] ), 
        .P2(\prop[0][3] ), .Gout(\gen[1][4] ), .Pout(\prop[1][4] ) );
  PG_53 PG1_2_1_3 ( .G1(\gen[0][6] ), .P1(\prop[0][6] ), .G2(\gen[0][5] ), 
        .P2(\prop[0][5] ), .Gout(\gen[1][6] ), .Pout(\prop[1][6] ) );
  PG_52 PG1_2_1_4 ( .G1(\gen[0][8] ), .P1(\prop[0][8] ), .G2(\gen[0][7] ), 
        .P2(\prop[0][7] ), .Gout(\gen[1][8] ), .Pout(\prop[1][8] ) );
  PG_51 PG1_2_1_5 ( .G1(\gen[0][10] ), .P1(\prop[0][10] ), .G2(\gen[0][9] ), 
        .P2(\prop[0][9] ), .Gout(\gen[1][10] ), .Pout(\prop[1][10] ) );
  PG_50 PG1_2_1_6 ( .G1(\gen[0][12] ), .P1(\prop[0][12] ), .G2(\gen[0][11] ), 
        .P2(\prop[0][11] ), .Gout(\gen[1][12] ), .Pout(\prop[1][12] ) );
  PG_49 PG1_2_1_7 ( .G1(\gen[0][14] ), .P1(\prop[0][14] ), .G2(\gen[0][13] ), 
        .P2(\prop[0][13] ), .Gout(\gen[1][14] ), .Pout(\prop[1][14] ) );
  PG_48 PG1_2_1_8 ( .G1(\gen[0][16] ), .P1(\prop[0][16] ), .G2(\gen[0][15] ), 
        .P2(\prop[0][15] ), .Gout(\gen[1][16] ), .Pout(\prop[1][16] ) );
  PG_47 PG1_2_1_9 ( .G1(\gen[0][18] ), .P1(\prop[0][18] ), .G2(\gen[0][17] ), 
        .P2(\prop[0][17] ), .Gout(\gen[1][18] ), .Pout(\prop[1][18] ) );
  PG_46 PG1_2_1_10 ( .G1(\gen[0][20] ), .P1(\prop[0][20] ), .G2(\gen[0][19] ), 
        .P2(\prop[0][19] ), .Gout(\gen[1][20] ), .Pout(\prop[1][20] ) );
  PG_45 PG1_2_1_11 ( .G1(\gen[0][22] ), .P1(\prop[0][22] ), .G2(\gen[0][21] ), 
        .P2(\prop[0][21] ), .Gout(\gen[1][22] ), .Pout(\prop[1][22] ) );
  PG_44 PG1_2_1_12 ( .G1(\gen[0][24] ), .P1(\prop[0][24] ), .G2(\gen[0][23] ), 
        .P2(\prop[0][23] ), .Gout(\gen[1][24] ), .Pout(\prop[1][24] ) );
  PG_43 PG1_2_1_13 ( .G1(\gen[0][26] ), .P1(\prop[0][26] ), .G2(\gen[0][25] ), 
        .P2(\prop[0][25] ), .Gout(\gen[1][26] ), .Pout(\prop[1][26] ) );
  PG_42 PG1_2_1_14 ( .G1(\gen[0][28] ), .P1(\prop[0][28] ), .G2(\gen[0][27] ), 
        .P2(\prop[0][27] ), .Gout(\gen[1][28] ), .Pout(\prop[1][28] ) );
  PG_41 PG1_2_1_15 ( .G1(\gen[0][30] ), .P1(\prop[0][30] ), .G2(\gen[0][29] ), 
        .P2(\prop[0][29] ), .Gout(\gen[1][30] ), .Pout(\prop[1][30] ) );
  PG_40 PG1_2_1_16 ( .G1(\gen[0][32] ), .P1(\prop[0][32] ), .G2(\gen[0][31] ), 
        .P2(\prop[0][31] ), .Gout(\gen[1][32] ), .Pout(\prop[1][32] ) );
  G_17 G1_2_2_1 ( .G1(\gen[1][4] ), .P1(\prop[1][4] ), .G2(\gen[1][2] ), 
        .Gout(n92) );
  PG_39 PG1_2_2_2 ( .G1(\gen[1][8] ), .P1(\prop[1][8] ), .G2(\gen[1][6] ), 
        .P2(\prop[1][6] ), .Gout(\gen[2][8] ), .Pout(\prop[2][8] ) );
  PG_38 PG1_2_2_3 ( .G1(\gen[1][12] ), .P1(\prop[1][12] ), .G2(\gen[1][10] ), 
        .P2(\prop[1][10] ), .Gout(n75), .Pout(\prop[2][12] ) );
  PG_37 PG1_2_2_4 ( .G1(\gen[1][16] ), .P1(\prop[1][16] ), .G2(\gen[1][14] ), 
        .P2(\prop[1][14] ), .Gout(\gen[2][16] ), .Pout(\prop[2][16] ) );
  PG_36 PG1_2_2_5 ( .G1(\gen[1][20] ), .P1(\prop[1][20] ), .G2(\gen[1][18] ), 
        .P2(\prop[1][18] ), .Gout(n79), .Pout(\prop[2][20] ) );
  PG_35 PG1_2_2_6 ( .G1(\gen[1][24] ), .P1(\prop[1][24] ), .G2(\gen[1][22] ), 
        .P2(\prop[1][22] ), .Gout(\gen[2][24] ), .Pout(\prop[2][24] ) );
  PG_34 PG1_2_2_7 ( .G1(\gen[1][28] ), .P1(\prop[1][28] ), .G2(\gen[1][26] ), 
        .P2(\prop[1][26] ), .Gout(n74), .Pout(\prop[2][28] ) );
  PG_33 PG1_2_2_8 ( .G1(\gen[1][32] ), .P1(\prop[1][32] ), .G2(\gen[1][30] ), 
        .P2(\prop[1][30] ), .Gout(\gen[2][32] ), .Pout(\prop[2][32] ) );
  G_16 G3_3_2 ( .G1(\gen[2][8] ), .P1(\prop[2][8] ), .G2(n92), .Gout(n81) );
  PG_32 PG3_3_4 ( .G1(\gen[2][16] ), .P1(\prop[2][16] ), .G2(n75), .P2(
        \prop[2][12] ), .Gout(\gen[3][16] ), .Pout(\prop[3][16] ) );
  PG_31 PG3_3_6 ( .G1(\gen[2][24] ), .P1(\prop[2][24] ), .G2(n79), .P2(
        \prop[2][20] ), .Gout(n78), .Pout(\prop[3][24] ) );
  PG_30 PG3_3_8 ( .G1(\gen[2][32] ), .P1(\prop[2][32] ), .G2(n74), .P2(
        \prop[2][28] ), .Gout(\gen[3][32] ), .Pout(\prop[3][32] ) );
  G_15 G3_E_4_2 ( .G1(n75), .P1(\prop[2][12] ), .G2(n89), .Gout(Cout[3]) );
  G_14 G3_E_4_3 ( .G1(\gen[3][16] ), .P1(\prop[3][16] ), .G2(n81), .Gout(n91)
         );
  PG_29 PG3_E_4_6 ( .G1(n74), .P1(\prop[2][28] ), .G2(n78), .P2(\prop[3][24] ), 
        .Gout(\gen[4][28] ), .Pout(\prop[4][28] ) );
  PG_28 PG3_E_4_7 ( .G1(\gen[3][32] ), .P1(\prop[3][32] ), .G2(n87), .P2(
        \prop[3][24] ), .Gout(\gen[4][32] ), .Pout(\prop[4][32] ) );
  G_13 G3_E_5_4 ( .G1(n86), .P1(\prop[2][20] ), .G2(n91), .Gout(Cout[5]) );
  G_12 G3_E_5_5 ( .G1(n87), .P1(\prop[3][24] ), .G2(n91), .Gout(Cout[6]) );
  G_11 G3_E_5_6 ( .G1(\gen[4][28] ), .P1(\prop[4][28] ), .G2(n91), .Gout(
        Cout[7]) );
  G_10 G3_E_5_7 ( .G1(\gen[4][32] ), .P1(\prop[4][32] ), .G2(Cout[4]), .Gout(
        Cout[8]) );
  BUF_X1 U1 ( .A(n89), .Z(Cout[2]) );
  BUF_X1 U2 ( .A(n92), .Z(Cout[1]) );
  CLKBUF_X1 U3 ( .A(n79), .Z(n86) );
  CLKBUF_X1 U4 ( .A(n78), .Z(n87) );
  BUF_X2 U5 ( .A(n91), .Z(Cout[4]) );
  CLKBUF_X1 U6 ( .A(n81), .Z(n89) );
  AOI21_X1 U7 ( .B1(propcin), .B2(Cin), .A(gencin), .ZN(n2) );
  INV_X1 U8 ( .A(n2), .ZN(\gen[0][1] ) );
endmodule


module BoothMulWallace_Nbit32_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29;

  XOR2_X1 U31 ( .A(A[9]), .B(n9), .Z(SUM[9]) );
  XOR2_X1 U32 ( .A(A[6]), .B(n12), .Z(SUM[6]) );
  XOR2_X1 U33 ( .A(A[4]), .B(n14), .Z(SUM[4]) );
  XOR2_X1 U34 ( .A(A[15]), .B(n19), .Z(SUM[15]) );
  XOR2_X1 U35 ( .A(A[13]), .B(n22), .Z(SUM[13]) );
  XOR2_X1 U36 ( .A(A[11]), .B(n25), .Z(SUM[11]) );
  NAND3_X1 U37 ( .A1(A[6]), .A2(n12), .A3(A[7]), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n17), .A2(n18), .ZN(n16) );
  NOR3_X1 U2 ( .A1(n18), .A2(n17), .A3(n15), .ZN(n14) );
  NOR2_X1 U3 ( .A1(n29), .A2(n13), .ZN(n12) );
  INV_X1 U4 ( .A(A[5]), .ZN(n29) );
  NOR2_X1 U5 ( .A1(n28), .A2(n10), .ZN(n9) );
  INV_X1 U6 ( .A(A[8]), .ZN(n28) );
  NOR2_X1 U7 ( .A1(n26), .A2(n27), .ZN(n25) );
  INV_X1 U8 ( .A(A[10]), .ZN(n26) );
  NOR2_X1 U9 ( .A1(n23), .A2(n24), .ZN(n22) );
  INV_X1 U10 ( .A(A[12]), .ZN(n23) );
  NAND2_X1 U11 ( .A1(A[1]), .A2(A[0]), .ZN(n17) );
  NAND2_X1 U12 ( .A1(n9), .A2(A[9]), .ZN(n27) );
  NAND2_X1 U13 ( .A1(A[4]), .A2(n14), .ZN(n13) );
  NAND2_X1 U14 ( .A1(A[11]), .A2(n25), .ZN(n24) );
  NAND2_X1 U15 ( .A1(A[13]), .A2(n22), .ZN(n20) );
  INV_X1 U16 ( .A(A[0]), .ZN(SUM[0]) );
  INV_X1 U17 ( .A(A[2]), .ZN(n18) );
  NAND2_X1 U18 ( .A1(A[6]), .A2(n12), .ZN(n11) );
  INV_X1 U19 ( .A(A[14]), .ZN(n21) );
  XNOR2_X1 U20 ( .A(A[14]), .B(n20), .ZN(SUM[14]) );
  XNOR2_X1 U21 ( .A(A[12]), .B(n24), .ZN(SUM[12]) );
  XNOR2_X1 U22 ( .A(A[8]), .B(n10), .ZN(SUM[8]) );
  XNOR2_X1 U23 ( .A(A[7]), .B(n11), .ZN(SUM[7]) );
  XNOR2_X1 U24 ( .A(n15), .B(n16), .ZN(SUM[3]) );
  XNOR2_X1 U25 ( .A(A[2]), .B(n17), .ZN(SUM[2]) );
  XNOR2_X1 U26 ( .A(A[5]), .B(n13), .ZN(SUM[5]) );
  XNOR2_X1 U27 ( .A(A[1]), .B(SUM[0]), .ZN(SUM[1]) );
  XNOR2_X1 U28 ( .A(A[10]), .B(n27), .ZN(SUM[10]) );
  NOR2_X1 U29 ( .A1(n20), .A2(n21), .ZN(n19) );
  INV_X1 U30 ( .A(A[3]), .ZN(n15) );
endmodule


module P4adderN_Nbit32 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;
  wire   n14, n7, n12, Carry_0_port, Carry_1_port, Carry_2_port, Carry_3_port,
         Carry_4_port, Carry_5_port, Carry_6_port, Carry_7_port, n9, n15, n21,
         n17, n16, n13, n20, n11, n18, n8, n2, n3, n5, n10, n1, n19, n6, n4;
  assign n14 = A[16];
  assign n7 = A[24];
  assign n12 = A[28];
  assign n9 = A[13];
  assign n15 = A[14];
  assign n21 = A[15];
  assign n17 = A[17];
  assign n16 = A[18];
  assign n13 = A[19];
  assign n20 = A[21];
  assign n11 = A[22];
  assign n18 = A[23];
  assign n8 = A[25];
  assign n2 = A[27];
  assign n3 = B[15];
  assign n5 = B[17];
  assign n10 = B[19];
  assign n1 = B[21];
  assign n19 = B[23];
  assign n6 = B[25];
  assign n4 = B[27];

  SparseTreeCarryGenNBM_Nbit32 STCG ( .A({A[31:29], n12, n2, A[26], n8, n7, 
        n18, n11, n20, A[20], n13, n16, n17, n14, n21, n15, n9, A[12:0]}), .B(
        {B[31:28], n4, B[26], n6, B[24], n19, B[22], n1, B[20], n10, B[18], n5, 
        B[16], n3, B[14:0]}), .Cin(Cin), .Cout({Cout, Carry_7_port, 
        Carry_6_port, Carry_5_port, Carry_4_port, Carry_3_port, Carry_2_port, 
        Carry_1_port, Carry_0_port}) );
  CarrySumNBM_Nbit32 CSN ( .A({A[31:29], n12, n2, A[26], n8, n7, n18, n11, n20, 
        A[20], n13, n16, n17, n14, n21, n15, n9, A[12:0]}), .B({B[31:28], n4, 
        B[26], n6, B[24], n19, B[22], n1, B[20], n10, B[18], n5, B[16], n3, 
        B[14:0]}), .Ci({Carry_7_port, Carry_6_port, Carry_5_port, Carry_4_port, 
        Carry_3_port, Carry_2_port, Carry_1_port, Carry_0_port}), .S(S) );
endmodule


module CSA_N32_1 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_96 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1]) );
  FA_95 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2]) );
  FA_94 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3]) );
  FA_93 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4]) );
  FA_92 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5]) );
  FA_91 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6]) );
  FA_90 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7]) );
  FA_89 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8]) );
  FA_88 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9]) );
  FA_87 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_86 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_85 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_84 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_83 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_82 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_81 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_80 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_79 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_78 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_77 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_76 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_75 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_74 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_73 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_72 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_71 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_70 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_69 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_68 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_67 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_66 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_65 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_2 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_128 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_127 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_126 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_125 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_124 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_123 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_122 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_121 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_120 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_119 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_118 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_117 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_116 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_115 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_114 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_113 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_112 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_111 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_110 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_109 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_108 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_107 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_106 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_105 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_104 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_103 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_102 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_101 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_100 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_99 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_98 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_97 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_3 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_160 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_159 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_158 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_157 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_156 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_155 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_154 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_153 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_152 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_151 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_150 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_149 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_148 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_147 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_146 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_145 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_144 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_143 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_142 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_141 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_140 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_139 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_138 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_137 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_136 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_135 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_134 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_133 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_132 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_131 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_130 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_129 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_4 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_192 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_191 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_190 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_189 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_188 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_187 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_186 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_185 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_184 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_183 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_182 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_181 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_180 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_179 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_178 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_177 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_176 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_175 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_174 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_173 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_172 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_171 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_170 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_169 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_168 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_167 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_166 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_165 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_164 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_163 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_162 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_161 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_5 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_224 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_223 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_222 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_221 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_220 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_219 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_218 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_217 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_216 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_215 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_214 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_213 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_212 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_211 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_210 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_209 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_208 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_207 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_206 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_205 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_204 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_203 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_202 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_201 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_200 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_199 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_198 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_197 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_196 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_195 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_194 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_193 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_6 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_256 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_255 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_254 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_253 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_252 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_251 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_250 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_249 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_248 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_247 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_246 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_245 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_244 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_243 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_242 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_241 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_240 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_239 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_238 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_237 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_236 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_235 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_234 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_233 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_232 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_231 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_230 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_229 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_228 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_227 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_226 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_225 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_7 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_288 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_287 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_286 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_285 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_284 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_283 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_282 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_281 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_280 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_279 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_278 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_277 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_276 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_275 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_274 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_273 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_272 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_271 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_270 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_269 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_268 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_267 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_266 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_265 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_264 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_263 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_262 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_261 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_260 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_259 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_258 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_257 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_8 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_320 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_319 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_318 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_317 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_316 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_315 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_314 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_313 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_312 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_311 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_310 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_309 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_308 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_307 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_306 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_305 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_304 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_303 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_302 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_301 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_300 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_299 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_298 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_297 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_296 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_295 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_294 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_293 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_292 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_291 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_290 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_289 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_9 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_352 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_351 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_350 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_349 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_348 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_347 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_346 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_345 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_344 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_343 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_342 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_341 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_340 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_339 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_338 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_337 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_336 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_335 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_334 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_333 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_332 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_331 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_330 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_329 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_328 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_327 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_326 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_325 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_324 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_323 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_322 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_321 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_10 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_384 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_383 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_382 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_381 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_380 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_379 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_378 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_377 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_376 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_375 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_374 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_373 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_372 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_371 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_370 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_369 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_368 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_367 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_366 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_365 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_364 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_363 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_362 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_361 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_360 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_359 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_358 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_357 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_356 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_355 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_354 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_353 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_11 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_416 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_415 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_414 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_413 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_412 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_411 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_410 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_409 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_408 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_407 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_406 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_405 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_404 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_403 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_402 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_401 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_400 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_399 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_398 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_397 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_396 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_395 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_394 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_393 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_392 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_391 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_390 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_389 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_388 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_387 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_386 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_385 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_12 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_448 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_447 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_446 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_445 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_444 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_443 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_442 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_441 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_440 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_439 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_438 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_437 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_436 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_435 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_434 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_433 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_432 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_431 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_430 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_429 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_428 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_427 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_426 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_425 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_424 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_423 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_422 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_421 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_420 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_419 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_418 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_417 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_13 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_480 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_479 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_478 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_477 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_476 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_475 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_474 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_473 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_472 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_471 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_470 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_469 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_468 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_467 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_466 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_465 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_464 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_463 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_462 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_461 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_460 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_459 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_458 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_457 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_456 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_455 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_454 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_453 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_452 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_451 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_450 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_449 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module CSA_N32_0 ( A, B, C, sum_out, cout );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  output [31:0] sum_out;
  output [31:0] cout;

  assign cout[0] = 1'b0;

  FA_0_0 st0_0 ( .A(A[0]), .B(B[0]), .Ci(C[0]), .S(sum_out[0]), .Co(cout[1])
         );
  FA_511 st0_1 ( .A(A[1]), .B(B[1]), .Ci(C[1]), .S(sum_out[1]), .Co(cout[2])
         );
  FA_510 st0_2 ( .A(A[2]), .B(B[2]), .Ci(C[2]), .S(sum_out[2]), .Co(cout[3])
         );
  FA_509 st0_3 ( .A(A[3]), .B(B[3]), .Ci(C[3]), .S(sum_out[3]), .Co(cout[4])
         );
  FA_508 st0_4 ( .A(A[4]), .B(B[4]), .Ci(C[4]), .S(sum_out[4]), .Co(cout[5])
         );
  FA_507 st0_5 ( .A(A[5]), .B(B[5]), .Ci(C[5]), .S(sum_out[5]), .Co(cout[6])
         );
  FA_506 st0_6 ( .A(A[6]), .B(B[6]), .Ci(C[6]), .S(sum_out[6]), .Co(cout[7])
         );
  FA_505 st0_7 ( .A(A[7]), .B(B[7]), .Ci(C[7]), .S(sum_out[7]), .Co(cout[8])
         );
  FA_504 st0_8 ( .A(A[8]), .B(B[8]), .Ci(C[8]), .S(sum_out[8]), .Co(cout[9])
         );
  FA_503 st0_9 ( .A(A[9]), .B(B[9]), .Ci(C[9]), .S(sum_out[9]), .Co(cout[10])
         );
  FA_502 st0_10 ( .A(A[10]), .B(B[10]), .Ci(C[10]), .S(sum_out[10]), .Co(
        cout[11]) );
  FA_501 st0_11 ( .A(A[11]), .B(B[11]), .Ci(C[11]), .S(sum_out[11]), .Co(
        cout[12]) );
  FA_500 st0_12 ( .A(A[12]), .B(B[12]), .Ci(C[12]), .S(sum_out[12]), .Co(
        cout[13]) );
  FA_499 st0_13 ( .A(A[13]), .B(B[13]), .Ci(C[13]), .S(sum_out[13]), .Co(
        cout[14]) );
  FA_498 st0_14 ( .A(A[14]), .B(B[14]), .Ci(C[14]), .S(sum_out[14]), .Co(
        cout[15]) );
  FA_497 st0_15 ( .A(A[15]), .B(B[15]), .Ci(C[15]), .S(sum_out[15]), .Co(
        cout[16]) );
  FA_496 st0_16 ( .A(A[16]), .B(B[16]), .Ci(C[16]), .S(sum_out[16]), .Co(
        cout[17]) );
  FA_495 st0_17 ( .A(A[17]), .B(B[17]), .Ci(C[17]), .S(sum_out[17]), .Co(
        cout[18]) );
  FA_494 st0_18 ( .A(A[18]), .B(B[18]), .Ci(C[18]), .S(sum_out[18]), .Co(
        cout[19]) );
  FA_493 st0_19 ( .A(A[19]), .B(B[19]), .Ci(C[19]), .S(sum_out[19]), .Co(
        cout[20]) );
  FA_492 st0_20 ( .A(A[20]), .B(B[20]), .Ci(C[20]), .S(sum_out[20]), .Co(
        cout[21]) );
  FA_491 st0_21 ( .A(A[21]), .B(B[21]), .Ci(C[21]), .S(sum_out[21]), .Co(
        cout[22]) );
  FA_490 st0_22 ( .A(A[22]), .B(B[22]), .Ci(C[22]), .S(sum_out[22]), .Co(
        cout[23]) );
  FA_489 st0_23 ( .A(A[23]), .B(B[23]), .Ci(C[23]), .S(sum_out[23]), .Co(
        cout[24]) );
  FA_488 st0_24 ( .A(A[24]), .B(B[24]), .Ci(C[24]), .S(sum_out[24]), .Co(
        cout[25]) );
  FA_487 st0_25 ( .A(A[25]), .B(B[25]), .Ci(C[25]), .S(sum_out[25]), .Co(
        cout[26]) );
  FA_486 st0_26 ( .A(A[26]), .B(B[26]), .Ci(C[26]), .S(sum_out[26]), .Co(
        cout[27]) );
  FA_485 st0_27 ( .A(A[27]), .B(B[27]), .Ci(C[27]), .S(sum_out[27]), .Co(
        cout[28]) );
  FA_484 st0_28 ( .A(A[28]), .B(B[28]), .Ci(C[28]), .S(sum_out[28]), .Co(
        cout[29]) );
  FA_483 st0_29 ( .A(A[29]), .B(B[29]), .Ci(C[29]), .S(sum_out[29]), .Co(
        cout[30]) );
  FA_482 st0_30 ( .A(A[30]), .B(B[30]), .Ci(C[30]), .S(sum_out[30]), .Co(
        cout[31]) );
  FA_481 st0_31 ( .A(A[31]), .B(B[31]), .Ci(C[31]), .S(sum_out[31]) );
endmodule


module MUX21_264 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_268 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_269 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_270 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_271 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_272 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_274 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_276 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_277 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_278 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_279 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_280 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_281 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_282 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_283 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_284 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_285 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_286 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_287 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_288 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_292 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n15;

  AOI22_X1 U1 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n15) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_294 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n16;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_296 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n18;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n18), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n18) );
endmodule


module MUX21_297 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n13;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n13) );
  AOI22_X1 U3 ( .A1(in0), .A2(n13), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_298 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n15;

  AOI22_X1 U1 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n15) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_299 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n14;

  INV_X1 U1 ( .A(S), .ZN(n14) );
  AOI22_X1 U2 ( .A1(in0), .A2(n14), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_300 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n13;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n13), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n13) );
endmodule


module MUX21_301 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n20;

  AOI22_X1 U1 ( .A1(n20), .A2(in0), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n20) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_302 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n14;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n14) );
  AOI22_X1 U3 ( .A1(in0), .A2(n14), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_303 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n12;

  AOI22_X1 U1 ( .A1(in0), .A2(n12), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n12) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_304 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n14;

  AOI22_X1 U1 ( .A1(in0), .A2(n14), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n14) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_305 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n15;

  INV_X1 U1 ( .A(S), .ZN(n15) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_306 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n14;

  AOI22_X1 U1 ( .A1(in0), .A2(n14), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n14) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_307 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n13;

  INV_X1 U1 ( .A(S), .ZN(n13) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n13), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_308 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n12;

  AOI22_X1 U1 ( .A1(in0), .A2(n12), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n12) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_309 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n9;

  INV_X1 U1 ( .A(S), .ZN(n9) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n9), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_310 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n17;

  INV_X1 U1 ( .A(S), .ZN(n17) );
  AOI22_X1 U2 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_311 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n9;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n9) );
  AOI22_X1 U3 ( .A1(in0), .A2(n9), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_312 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n10;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n10) );
endmodule


module MUX21_313 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n21;

  INV_X1 U1 ( .A(S), .ZN(n21) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n21), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_314 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n21;

  AOI22_X1 U1 ( .A1(in0), .A2(n21), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n21) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_315 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n10;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n10) );
  AOI22_X1 U3 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_316 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n13;

  INV_X1 U1 ( .A(S), .ZN(n13) );
  AOI22_X1 U2 ( .A1(in0), .A2(n13), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_317 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n16;

  INV_X1 U1 ( .A(S), .ZN(n16) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n16), .A2(in0), .B1(S), .B2(in1), .ZN(n3) );
endmodule


module MUX21_318 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n13;

  INV_X1 U1 ( .A(S), .ZN(n13) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n13), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_319 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n13;

  INV_X1 U1 ( .A(S), .ZN(n13) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n13), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_320 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n8;

  INV_X1 U1 ( .A(S), .ZN(n8) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n8), .B1(S), .B2(in1), .ZN(n3) );
endmodule


module MUX21_322 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n12;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n12), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n12) );
endmodule


module MUX21_323 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n9;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n9), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n9) );
endmodule


module MUX21_324 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n10;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n10) );
endmodule


module MUX21_327 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n15;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n15) );
endmodule


module MUX21_328 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n14;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n14), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n14) );
endmodule


module MUX21_329 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n10;

  AOI22_X1 U1 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n10) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_330 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n14;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n14), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n14) );
endmodule


module MUX21_331 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n16;

  AOI22_X1 U1 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n16) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_332 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n15;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n15) );
endmodule


module MUX21_333 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n11;

  AOI22_X1 U1 ( .A1(in0), .A2(n11), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n11) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_334 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n14;

  AOI22_X1 U1 ( .A1(in0), .A2(n14), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n14) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_335 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n12;

  AOI22_X1 U1 ( .A1(in0), .A2(n12), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n12) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_336 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n12;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n12), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n12) );
endmodule


module MUX21_337 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n8;

  INV_X1 U1 ( .A(S), .ZN(n8) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n8), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_338 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n14;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  INV_X1 U2 ( .A(S), .ZN(n14) );
  AOI22_X1 U3 ( .A1(in0), .A2(n14), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_339 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n10;

  INV_X1 U1 ( .A(S), .ZN(n10) );
  AOI22_X1 U2 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_340 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n19;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n19), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n19) );
endmodule


module MUX21_341 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n15;

  INV_X1 U1 ( .A(S), .ZN(n15) );
  AOI22_X1 U2 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_342 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n9;

  AOI22_X1 U1 ( .A1(in0), .A2(n9), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n9) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_343 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n11;

  INV_X1 U1 ( .A(S), .ZN(n11) );
  AOI22_X1 U2 ( .A1(in0), .A2(n11), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_344 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n13;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n13), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n13) );
endmodule


module MUX21_345 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n12;

  INV_X1 U1 ( .A(S), .ZN(n12) );
  AOI22_X1 U2 ( .A1(in0), .A2(n12), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_346 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n17;

  AOI22_X1 U1 ( .A1(in0), .A2(n17), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n17) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_347 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n10;

  AOI22_X1 U1 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n10) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_348 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n10;

  AOI22_X1 U1 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n10) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_349 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n8;

  INV_X1 U1 ( .A(S), .ZN(n8) );
  AOI22_X1 U2 ( .A1(in0), .A2(n8), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_350 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n10;

  INV_X1 U1 ( .A(S), .ZN(n10) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_351 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n19;

  AOI22_X1 U1 ( .A1(in0), .A2(n19), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n19) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_352 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n5;

  INV_X1 U1 ( .A(S), .ZN(n5) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n5), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module CSBlockN_Nbit4_9 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_34 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_33 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_17 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_10 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_36 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_35 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_18 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_11 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_38 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_37 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_19 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_12 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_40 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_39 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_20 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_13 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_42 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_41 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_21 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_14 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_44 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_43 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_22 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_15 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_46 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_45 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_23 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_16 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_48 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_47 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_24 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module PG_55 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module G_27 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module MUX21_363 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_364 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_365 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_366 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_367 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module CSBlockN_Nbit4_17 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_50 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_49 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_25 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_18 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_52 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_51 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_26 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_19 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_54 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_53 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_27 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_20 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_56 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_55 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_28 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_21 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_58 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_57 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_29 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_22 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_60 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_59 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_30 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_23 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_62 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_61 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_31 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module CSBlockN_Nbit4_0 ( A, B, Ci, S, Cout );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Cout;

  wire   [4:0] sum_cin0;
  wire   [4:0] sum_cin1;

  RCAN_Nbit4_16 RCA_Cin_0 ( .A(A), .B(B), .Ci(1'b0), .S(sum_cin0[3:0]), .Co(
        sum_cin0[4]) );
  RCAN_Nbit4_63 RCA_Cin_1 ( .A(A), .B(B), .Ci(1'b1), .S(sum_cin1[3:0]), .Co(
        sum_cin1[4]) );
  mux21N_N5_32 MUX ( .in1(sum_cin1), .in0(sum_cin0), .S(Ci), .U({Cout, S}) );
endmodule


module G_28 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_29 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_30 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_31 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PG_82 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P2), .A2(P1), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module G_32 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module G_33 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PG_86 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module G_34 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PG_93 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module G_35 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PG_94 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_95 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_98 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_99 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_100 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_101 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_102 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module PG_103 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_104 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_105 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_106 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_107 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P2), .A2(P1), .ZN(Pout) );
endmodule


module PG_27 ( G1, P1, G2, P2, Gout, Pout );
  input G1, P1, G2, P2;
  output Gout, Pout;
  wire   n2;

  AND2_X1 U1 ( .A1(P2), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G2), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module G_9 ( G1, P1, G2, Gout );
  input G1, P1, G2;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G2), .A(G1), .ZN(n2) );
endmodule


module PGblock_121 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_122 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_123 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_124 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_125 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_126 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_127 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGblock_32 ( A, B, G, P );
  input A, B;
  output G, P;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module mux21N_N32_1 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;


  MUX21_192 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_191 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_190 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_189 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_188 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
  MUX21_187 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(S), .Y(U[5]) );
  MUX21_186 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(S), .Y(U[6]) );
  MUX21_185 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(S), .Y(U[7]) );
  MUX21_184 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(S), .Y(U[8]) );
  MUX21_183 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(S), .Y(U[9]) );
  MUX21_182 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(S), .Y(U[10]) );
  MUX21_181 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(S), .Y(U[11]) );
  MUX21_180 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(S), .Y(U[12]) );
  MUX21_179 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(S), .Y(U[13]) );
  MUX21_178 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(S), .Y(U[14]) );
  MUX21_177 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(S), .Y(U[15]) );
  MUX21_176 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(S), .Y(U[16]) );
  MUX21_175 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(S), .Y(U[17]) );
  MUX21_174 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(S), .Y(U[18]) );
  MUX21_173 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(S), .Y(U[19]) );
  MUX21_172 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(S), .Y(U[20]) );
  MUX21_171 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(S), .Y(U[21]) );
  MUX21_170 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(S), .Y(U[22]) );
  MUX21_169 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(S), .Y(U[23]) );
  MUX21_168 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(S), .Y(U[24]) );
  MUX21_167 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(S), .Y(U[25]) );
  MUX21_166 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(S), .Y(U[26]) );
  MUX21_165 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(S), .Y(U[27]) );
  MUX21_164 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(S), .Y(U[28]) );
  MUX21_163 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(S), .Y(U[29]) );
  MUX21_162 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(S), .Y(U[30]) );
  MUX21_161 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(S), .Y(U[31]) );
endmodule


module mux21N_N32_2 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;


  MUX21_224 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_223 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_222 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_221 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_220 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
  MUX21_219 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(S), .Y(U[5]) );
  MUX21_218 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(S), .Y(U[6]) );
  MUX21_217 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(S), .Y(U[7]) );
  MUX21_216 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(S), .Y(U[8]) );
  MUX21_215 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(S), .Y(U[9]) );
  MUX21_214 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(S), .Y(U[10]) );
  MUX21_213 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(S), .Y(U[11]) );
  MUX21_212 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(S), .Y(U[12]) );
  MUX21_211 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(S), .Y(U[13]) );
  MUX21_210 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(S), .Y(U[14]) );
  MUX21_209 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(S), .Y(U[15]) );
  MUX21_208 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(S), .Y(U[16]) );
  MUX21_207 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(S), .Y(U[17]) );
  MUX21_206 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(S), .Y(U[18]) );
  MUX21_205 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(S), .Y(U[19]) );
  MUX21_204 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(S), .Y(U[20]) );
  MUX21_203 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(S), .Y(U[21]) );
  MUX21_202 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(S), .Y(U[22]) );
  MUX21_201 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(S), .Y(U[23]) );
  MUX21_200 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(S), .Y(U[24]) );
  MUX21_199 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(S), .Y(U[25]) );
  MUX21_198 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(S), .Y(U[26]) );
  MUX21_197 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(S), .Y(U[27]) );
  MUX21_196 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(S), .Y(U[28]) );
  MUX21_195 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(S), .Y(U[29]) );
  MUX21_194 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(S), .Y(U[30]) );
  MUX21_193 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(S), .Y(U[31]) );
endmodule


module mux21N_N32_3 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;


  MUX21_256 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_255 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_254 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_253 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_252 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
  MUX21_251 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(S), .Y(U[5]) );
  MUX21_250 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(S), .Y(U[6]) );
  MUX21_249 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(S), .Y(U[7]) );
  MUX21_248 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(S), .Y(U[8]) );
  MUX21_247 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(S), .Y(U[9]) );
  MUX21_246 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(S), .Y(U[10]) );
  MUX21_245 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(S), .Y(U[11]) );
  MUX21_244 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(S), .Y(U[12]) );
  MUX21_243 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(S), .Y(U[13]) );
  MUX21_242 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(S), .Y(U[14]) );
  MUX21_241 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(S), .Y(U[15]) );
  MUX21_240 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(S), .Y(U[16]) );
  MUX21_239 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(S), .Y(U[17]) );
  MUX21_238 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(S), .Y(U[18]) );
  MUX21_237 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(S), .Y(U[19]) );
  MUX21_236 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(S), .Y(U[20]) );
  MUX21_235 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(S), .Y(U[21]) );
  MUX21_234 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(S), .Y(U[22]) );
  MUX21_233 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(S), .Y(U[23]) );
  MUX21_232 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(S), .Y(U[24]) );
  MUX21_231 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(S), .Y(U[25]) );
  MUX21_230 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(S), .Y(U[26]) );
  MUX21_229 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(S), .Y(U[27]) );
  MUX21_228 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(S), .Y(U[28]) );
  MUX21_227 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(S), .Y(U[29]) );
  MUX21_226 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(S), .Y(U[30]) );
  MUX21_225 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(S), .Y(U[31]) );
endmodule


module MUX21_432 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_434 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  AOI22_X1 U1 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U2 ( .A(S), .ZN(n4) );
  INV_X1 U3 ( .A(n3), .ZN(Y) );
endmodule


module MUX21_435 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_436 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_437 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_438 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module LogicFun_v2_Nbit32 ( A, B, notA, notB, AandB, AorB, AxorB, AnandB, 
        AnorB, AxnorB );
  input [31:0] A;
  input [31:0] B;
  output [31:0] notA;
  output [31:0] notB;
  output [31:0] AandB;
  output [31:0] AorB;
  output [31:0] AxorB;
  output [31:0] AnandB;
  output [31:0] AnorB;
  output [31:0] AxnorB;


  INV_X1 U1 ( .A(AxorB[1]), .ZN(AxnorB[1]) );
  INV_X1 U2 ( .A(AxorB[0]), .ZN(AxnorB[0]) );
  INV_X1 U3 ( .A(AxorB[15]), .ZN(AxnorB[15]) );
  INV_X1 U4 ( .A(AxorB[10]), .ZN(AxnorB[10]) );
  INV_X1 U5 ( .A(AxorB[11]), .ZN(AxnorB[11]) );
  INV_X1 U6 ( .A(AxorB[12]), .ZN(AxnorB[12]) );
  INV_X1 U7 ( .A(AxorB[16]), .ZN(AxnorB[16]) );
  INV_X1 U8 ( .A(AxorB[17]), .ZN(AxnorB[17]) );
  INV_X1 U9 ( .A(AxorB[18]), .ZN(AxnorB[18]) );
  INV_X1 U10 ( .A(AxorB[23]), .ZN(AxnorB[23]) );
  INV_X1 U11 ( .A(AxorB[24]), .ZN(AxnorB[24]) );
  INV_X1 U12 ( .A(AxorB[25]), .ZN(AxnorB[25]) );
  INV_X1 U13 ( .A(AxorB[29]), .ZN(AxnorB[29]) );
  INV_X1 U14 ( .A(AxorB[30]), .ZN(AxnorB[30]) );
  INV_X1 U15 ( .A(AxorB[5]), .ZN(AxnorB[5]) );
  XNOR2_X1 U16 ( .A(notA[1]), .B(B[1]), .ZN(AxorB[1]) );
  XNOR2_X1 U17 ( .A(notA[0]), .B(B[0]), .ZN(AxorB[0]) );
  XNOR2_X1 U18 ( .A(notA[15]), .B(B[15]), .ZN(AxorB[15]) );
  XNOR2_X1 U19 ( .A(notA[10]), .B(B[10]), .ZN(AxorB[10]) );
  XNOR2_X1 U20 ( .A(notA[12]), .B(B[12]), .ZN(AxorB[12]) );
  XNOR2_X1 U21 ( .A(notA[11]), .B(B[11]), .ZN(AxorB[11]) );
  XNOR2_X1 U22 ( .A(notA[16]), .B(B[16]), .ZN(AxorB[16]) );
  XNOR2_X1 U23 ( .A(notA[17]), .B(B[17]), .ZN(AxorB[17]) );
  XNOR2_X1 U24 ( .A(notA[18]), .B(B[18]), .ZN(AxorB[18]) );
  XNOR2_X1 U25 ( .A(notA[23]), .B(B[23]), .ZN(AxorB[23]) );
  XNOR2_X1 U26 ( .A(notA[24]), .B(B[24]), .ZN(AxorB[24]) );
  XNOR2_X1 U27 ( .A(notA[25]), .B(B[25]), .ZN(AxorB[25]) );
  XNOR2_X1 U28 ( .A(notA[29]), .B(B[29]), .ZN(AxorB[29]) );
  XNOR2_X1 U29 ( .A(notA[30]), .B(B[30]), .ZN(AxorB[30]) );
  XNOR2_X1 U30 ( .A(notA[5]), .B(B[5]), .ZN(AxorB[5]) );
  INV_X1 U31 ( .A(B[1]), .ZN(notB[1]) );
  INV_X1 U32 ( .A(B[15]), .ZN(notB[15]) );
  INV_X1 U33 ( .A(B[0]), .ZN(notB[0]) );
  INV_X1 U34 ( .A(B[24]), .ZN(notB[24]) );
  INV_X1 U35 ( .A(B[23]), .ZN(notB[23]) );
  INV_X1 U36 ( .A(B[18]), .ZN(notB[18]) );
  INV_X1 U37 ( .A(B[17]), .ZN(notB[17]) );
  INV_X1 U38 ( .A(B[16]), .ZN(notB[16]) );
  INV_X1 U39 ( .A(B[29]), .ZN(notB[29]) );
  INV_X1 U40 ( .A(B[25]), .ZN(notB[25]) );
  INV_X1 U41 ( .A(B[30]), .ZN(notB[30]) );
  INV_X1 U42 ( .A(B[12]), .ZN(notB[12]) );
  INV_X1 U43 ( .A(B[10]), .ZN(notB[10]) );
  INV_X1 U44 ( .A(B[11]), .ZN(notB[11]) );
  INV_X1 U45 ( .A(B[5]), .ZN(notB[5]) );
  INV_X1 U46 ( .A(AxorB[19]), .ZN(AxnorB[19]) );
  INV_X1 U47 ( .A(AxorB[14]), .ZN(AxnorB[14]) );
  INV_X1 U48 ( .A(AxorB[13]), .ZN(AxnorB[13]) );
  INV_X1 U49 ( .A(AxorB[2]), .ZN(AxnorB[2]) );
  INV_X1 U50 ( .A(AxorB[3]), .ZN(AxnorB[3]) );
  INV_X1 U51 ( .A(AxorB[8]), .ZN(AxnorB[8]) );
  INV_X1 U52 ( .A(AxorB[20]), .ZN(AxnorB[20]) );
  INV_X1 U53 ( .A(AxorB[21]), .ZN(AxnorB[21]) );
  INV_X1 U54 ( .A(AxorB[22]), .ZN(AxnorB[22]) );
  INV_X1 U55 ( .A(AxorB[26]), .ZN(AxnorB[26]) );
  INV_X1 U56 ( .A(AxorB[27]), .ZN(AxnorB[27]) );
  INV_X1 U57 ( .A(AxorB[28]), .ZN(AxnorB[28]) );
  INV_X1 U58 ( .A(AxorB[31]), .ZN(AxnorB[31]) );
  INV_X1 U59 ( .A(AxorB[4]), .ZN(AxnorB[4]) );
  INV_X1 U60 ( .A(AxorB[6]), .ZN(AxnorB[6]) );
  INV_X1 U61 ( .A(AxorB[7]), .ZN(AxnorB[7]) );
  INV_X1 U62 ( .A(AxorB[9]), .ZN(AxnorB[9]) );
  INV_X1 U63 ( .A(AorB[25]), .ZN(AnorB[25]) );
  NAND2_X1 U64 ( .A1(notB[25]), .A2(notA[25]), .ZN(AorB[25]) );
  INV_X1 U65 ( .A(AorB[31]), .ZN(AnorB[31]) );
  NAND2_X1 U66 ( .A1(notB[31]), .A2(notA[31]), .ZN(AorB[31]) );
  INV_X1 U67 ( .A(AorB[29]), .ZN(AnorB[29]) );
  NAND2_X1 U68 ( .A1(notB[29]), .A2(notA[29]), .ZN(AorB[29]) );
  INV_X1 U69 ( .A(AorB[28]), .ZN(AnorB[28]) );
  NAND2_X1 U70 ( .A1(notB[28]), .A2(notA[28]), .ZN(AorB[28]) );
  XNOR2_X1 U71 ( .A(notA[14]), .B(B[14]), .ZN(AxorB[14]) );
  XNOR2_X1 U72 ( .A(notA[19]), .B(B[19]), .ZN(AxorB[19]) );
  XNOR2_X1 U73 ( .A(notA[13]), .B(B[13]), .ZN(AxorB[13]) );
  XNOR2_X1 U74 ( .A(notA[2]), .B(B[2]), .ZN(AxorB[2]) );
  XNOR2_X1 U75 ( .A(notA[3]), .B(B[3]), .ZN(AxorB[3]) );
  XNOR2_X1 U76 ( .A(notA[8]), .B(B[8]), .ZN(AxorB[8]) );
  XNOR2_X1 U77 ( .A(notA[20]), .B(B[20]), .ZN(AxorB[20]) );
  XNOR2_X1 U78 ( .A(notA[21]), .B(B[21]), .ZN(AxorB[21]) );
  XNOR2_X1 U79 ( .A(notA[22]), .B(B[22]), .ZN(AxorB[22]) );
  XNOR2_X1 U80 ( .A(notA[26]), .B(B[26]), .ZN(AxorB[26]) );
  XNOR2_X1 U81 ( .A(notA[27]), .B(B[27]), .ZN(AxorB[27]) );
  XNOR2_X1 U82 ( .A(notA[28]), .B(B[28]), .ZN(AxorB[28]) );
  XNOR2_X1 U83 ( .A(notA[31]), .B(B[31]), .ZN(AxorB[31]) );
  XNOR2_X1 U84 ( .A(notA[4]), .B(B[4]), .ZN(AxorB[4]) );
  XNOR2_X1 U85 ( .A(notA[6]), .B(B[6]), .ZN(AxorB[6]) );
  XNOR2_X1 U86 ( .A(notA[7]), .B(B[7]), .ZN(AxorB[7]) );
  XNOR2_X1 U87 ( .A(notA[9]), .B(B[9]), .ZN(AxorB[9]) );
  INV_X1 U88 ( .A(AorB[27]), .ZN(AnorB[27]) );
  NAND2_X1 U89 ( .A1(notB[27]), .A2(notA[27]), .ZN(AorB[27]) );
  INV_X1 U90 ( .A(AorB[26]), .ZN(AnorB[26]) );
  NAND2_X1 U91 ( .A1(notB[26]), .A2(notA[26]), .ZN(AorB[26]) );
  INV_X1 U92 ( .A(AorB[24]), .ZN(AnorB[24]) );
  NAND2_X1 U93 ( .A1(notB[24]), .A2(notA[24]), .ZN(AorB[24]) );
  INV_X1 U94 ( .A(AorB[23]), .ZN(AnorB[23]) );
  NAND2_X1 U95 ( .A1(notB[23]), .A2(notA[23]), .ZN(AorB[23]) );
  INV_X1 U96 ( .A(AorB[22]), .ZN(AnorB[22]) );
  NAND2_X1 U97 ( .A1(notB[22]), .A2(notA[22]), .ZN(AorB[22]) );
  INV_X1 U98 ( .A(AorB[21]), .ZN(AnorB[21]) );
  NAND2_X1 U99 ( .A1(notB[21]), .A2(notA[21]), .ZN(AorB[21]) );
  INV_X1 U100 ( .A(AorB[20]), .ZN(AnorB[20]) );
  NAND2_X1 U101 ( .A1(notB[20]), .A2(notA[20]), .ZN(AorB[20]) );
  INV_X1 U102 ( .A(AorB[30]), .ZN(AnorB[30]) );
  NAND2_X1 U103 ( .A1(notB[30]), .A2(notA[30]), .ZN(AorB[30]) );
  INV_X1 U104 ( .A(AorB[19]), .ZN(AnorB[19]) );
  NAND2_X1 U105 ( .A1(notB[19]), .A2(notA[19]), .ZN(AorB[19]) );
  INV_X1 U106 ( .A(AorB[18]), .ZN(AnorB[18]) );
  NAND2_X1 U107 ( .A1(notB[18]), .A2(notA[18]), .ZN(AorB[18]) );
  INV_X1 U108 ( .A(AorB[17]), .ZN(AnorB[17]) );
  NAND2_X1 U109 ( .A1(notB[17]), .A2(notA[17]), .ZN(AorB[17]) );
  INV_X1 U110 ( .A(AorB[16]), .ZN(AnorB[16]) );
  NAND2_X1 U111 ( .A1(notB[16]), .A2(notA[16]), .ZN(AorB[16]) );
  INV_X1 U112 ( .A(AorB[15]), .ZN(AnorB[15]) );
  NAND2_X1 U113 ( .A1(notB[15]), .A2(notA[15]), .ZN(AorB[15]) );
  INV_X1 U114 ( .A(AorB[14]), .ZN(AnorB[14]) );
  NAND2_X1 U115 ( .A1(notB[14]), .A2(notA[14]), .ZN(AorB[14]) );
  INV_X1 U116 ( .A(AorB[13]), .ZN(AnorB[13]) );
  NAND2_X1 U117 ( .A1(notB[13]), .A2(notA[13]), .ZN(AorB[13]) );
  INV_X1 U118 ( .A(AorB[12]), .ZN(AnorB[12]) );
  NAND2_X1 U119 ( .A1(notB[12]), .A2(notA[12]), .ZN(AorB[12]) );
  INV_X1 U120 ( .A(AorB[11]), .ZN(AnorB[11]) );
  NAND2_X1 U121 ( .A1(notB[11]), .A2(notA[11]), .ZN(AorB[11]) );
  INV_X1 U122 ( .A(AorB[10]), .ZN(AnorB[10]) );
  NAND2_X1 U123 ( .A1(notB[10]), .A2(notA[10]), .ZN(AorB[10]) );
  INV_X1 U124 ( .A(AorB[9]), .ZN(AnorB[9]) );
  NAND2_X1 U125 ( .A1(notB[9]), .A2(notA[9]), .ZN(AorB[9]) );
  INV_X1 U126 ( .A(AorB[8]), .ZN(AnorB[8]) );
  NAND2_X1 U127 ( .A1(notB[8]), .A2(notA[8]), .ZN(AorB[8]) );
  INV_X1 U128 ( .A(AorB[7]), .ZN(AnorB[7]) );
  NAND2_X1 U129 ( .A1(notB[7]), .A2(notA[7]), .ZN(AorB[7]) );
  INV_X1 U130 ( .A(AorB[6]), .ZN(AnorB[6]) );
  NAND2_X1 U131 ( .A1(notB[6]), .A2(notA[6]), .ZN(AorB[6]) );
  INV_X1 U132 ( .A(AorB[5]), .ZN(AnorB[5]) );
  NAND2_X1 U133 ( .A1(notB[5]), .A2(notA[5]), .ZN(AorB[5]) );
  INV_X1 U134 ( .A(AorB[4]), .ZN(AnorB[4]) );
  NAND2_X1 U135 ( .A1(notB[4]), .A2(notA[4]), .ZN(AorB[4]) );
  INV_X1 U136 ( .A(AorB[3]), .ZN(AnorB[3]) );
  NAND2_X1 U137 ( .A1(notB[3]), .A2(notA[3]), .ZN(AorB[3]) );
  INV_X1 U138 ( .A(AorB[2]), .ZN(AnorB[2]) );
  NAND2_X1 U139 ( .A1(notB[2]), .A2(notA[2]), .ZN(AorB[2]) );
  INV_X1 U140 ( .A(AorB[1]), .ZN(AnorB[1]) );
  NAND2_X1 U141 ( .A1(notB[1]), .A2(notA[1]), .ZN(AorB[1]) );
  INV_X1 U142 ( .A(AorB[0]), .ZN(AnorB[0]) );
  NAND2_X1 U143 ( .A1(notB[0]), .A2(notA[0]), .ZN(AorB[0]) );
  INV_X1 U144 ( .A(B[19]), .ZN(notB[19]) );
  INV_X1 U145 ( .A(B[14]), .ZN(notB[14]) );
  INV_X1 U146 ( .A(B[13]), .ZN(notB[13]) );
  INV_X1 U147 ( .A(B[8]), .ZN(notB[8]) );
  INV_X1 U148 ( .A(B[3]), .ZN(notB[3]) );
  INV_X1 U149 ( .A(B[2]), .ZN(notB[2]) );
  INV_X1 U150 ( .A(A[31]), .ZN(notA[31]) );
  INV_X1 U151 ( .A(A[30]), .ZN(notA[30]) );
  INV_X1 U152 ( .A(A[29]), .ZN(notA[29]) );
  INV_X1 U153 ( .A(A[28]), .ZN(notA[28]) );
  INV_X1 U154 ( .A(A[27]), .ZN(notA[27]) );
  INV_X1 U155 ( .A(A[26]), .ZN(notA[26]) );
  INV_X1 U156 ( .A(A[25]), .ZN(notA[25]) );
  INV_X1 U157 ( .A(A[24]), .ZN(notA[24]) );
  INV_X1 U158 ( .A(A[23]), .ZN(notA[23]) );
  INV_X1 U159 ( .A(A[22]), .ZN(notA[22]) );
  INV_X1 U160 ( .A(A[21]), .ZN(notA[21]) );
  INV_X1 U161 ( .A(A[20]), .ZN(notA[20]) );
  INV_X1 U162 ( .A(A[19]), .ZN(notA[19]) );
  INV_X1 U163 ( .A(A[18]), .ZN(notA[18]) );
  INV_X1 U164 ( .A(A[17]), .ZN(notA[17]) );
  INV_X1 U165 ( .A(A[16]), .ZN(notA[16]) );
  INV_X1 U166 ( .A(A[15]), .ZN(notA[15]) );
  INV_X1 U167 ( .A(A[14]), .ZN(notA[14]) );
  INV_X1 U168 ( .A(A[6]), .ZN(notA[6]) );
  INV_X1 U169 ( .A(A[5]), .ZN(notA[5]) );
  INV_X1 U170 ( .A(A[4]), .ZN(notA[4]) );
  INV_X1 U171 ( .A(A[3]), .ZN(notA[3]) );
  INV_X1 U172 ( .A(A[2]), .ZN(notA[2]) );
  INV_X1 U173 ( .A(A[1]), .ZN(notA[1]) );
  INV_X1 U174 ( .A(A[13]), .ZN(notA[13]) );
  INV_X1 U175 ( .A(A[12]), .ZN(notA[12]) );
  INV_X1 U176 ( .A(A[11]), .ZN(notA[11]) );
  INV_X1 U177 ( .A(A[10]), .ZN(notA[10]) );
  INV_X1 U178 ( .A(A[9]), .ZN(notA[9]) );
  INV_X1 U179 ( .A(A[8]), .ZN(notA[8]) );
  INV_X1 U180 ( .A(A[7]), .ZN(notA[7]) );
  INV_X1 U181 ( .A(A[0]), .ZN(notA[0]) );
  INV_X1 U182 ( .A(B[26]), .ZN(notB[26]) );
  INV_X1 U183 ( .A(B[22]), .ZN(notB[22]) );
  INV_X1 U184 ( .A(B[20]), .ZN(notB[20]) );
  INV_X1 U185 ( .A(B[31]), .ZN(notB[31]) );
  INV_X1 U186 ( .A(B[28]), .ZN(notB[28]) );
  INV_X1 U187 ( .A(B[27]), .ZN(notB[27]) );
  INV_X1 U188 ( .A(B[21]), .ZN(notB[21]) );
  INV_X1 U189 ( .A(B[9]), .ZN(notB[9]) );
  INV_X1 U190 ( .A(B[7]), .ZN(notB[7]) );
  INV_X1 U191 ( .A(B[6]), .ZN(notB[6]) );
  INV_X1 U192 ( .A(B[4]), .ZN(notB[4]) );
  INV_X1 U193 ( .A(AnandB[19]), .ZN(AandB[19]) );
  NAND2_X1 U194 ( .A1(A[19]), .A2(B[19]), .ZN(AnandB[19]) );
  INV_X1 U195 ( .A(AnandB[15]), .ZN(AandB[15]) );
  NAND2_X1 U196 ( .A1(A[15]), .A2(B[15]), .ZN(AnandB[15]) );
  INV_X1 U197 ( .A(AnandB[14]), .ZN(AandB[14]) );
  NAND2_X1 U198 ( .A1(A[14]), .A2(B[14]), .ZN(AnandB[14]) );
  INV_X1 U199 ( .A(AnandB[13]), .ZN(AandB[13]) );
  NAND2_X1 U200 ( .A1(A[13]), .A2(B[13]), .ZN(AnandB[13]) );
  INV_X1 U201 ( .A(AnandB[8]), .ZN(AandB[8]) );
  NAND2_X1 U202 ( .A1(A[8]), .A2(B[8]), .ZN(AnandB[8]) );
  INV_X1 U203 ( .A(AnandB[3]), .ZN(AandB[3]) );
  NAND2_X1 U204 ( .A1(A[3]), .A2(B[3]), .ZN(AnandB[3]) );
  INV_X1 U205 ( .A(AnandB[2]), .ZN(AandB[2]) );
  NAND2_X1 U206 ( .A1(A[2]), .A2(B[2]), .ZN(AnandB[2]) );
  INV_X1 U207 ( .A(AnandB[1]), .ZN(AandB[1]) );
  NAND2_X1 U208 ( .A1(A[1]), .A2(B[1]), .ZN(AnandB[1]) );
  INV_X1 U209 ( .A(AnandB[0]), .ZN(AandB[0]) );
  NAND2_X1 U210 ( .A1(A[0]), .A2(B[0]), .ZN(AnandB[0]) );
  INV_X1 U211 ( .A(AnandB[31]), .ZN(AandB[31]) );
  NAND2_X1 U212 ( .A1(A[31]), .A2(B[31]), .ZN(AnandB[31]) );
  INV_X1 U213 ( .A(AnandB[30]), .ZN(AandB[30]) );
  NAND2_X1 U214 ( .A1(A[30]), .A2(B[30]), .ZN(AnandB[30]) );
  INV_X1 U215 ( .A(AnandB[29]), .ZN(AandB[29]) );
  NAND2_X1 U216 ( .A1(A[29]), .A2(B[29]), .ZN(AnandB[29]) );
  INV_X1 U217 ( .A(AnandB[28]), .ZN(AandB[28]) );
  NAND2_X1 U218 ( .A1(A[28]), .A2(B[28]), .ZN(AnandB[28]) );
  INV_X1 U219 ( .A(AnandB[27]), .ZN(AandB[27]) );
  NAND2_X1 U220 ( .A1(A[27]), .A2(B[27]), .ZN(AnandB[27]) );
  INV_X1 U221 ( .A(AnandB[26]), .ZN(AandB[26]) );
  NAND2_X1 U222 ( .A1(A[26]), .A2(B[26]), .ZN(AnandB[26]) );
  INV_X1 U223 ( .A(AnandB[25]), .ZN(AandB[25]) );
  NAND2_X1 U224 ( .A1(A[25]), .A2(B[25]), .ZN(AnandB[25]) );
  INV_X1 U225 ( .A(AnandB[24]), .ZN(AandB[24]) );
  NAND2_X1 U226 ( .A1(A[24]), .A2(B[24]), .ZN(AnandB[24]) );
  INV_X1 U227 ( .A(AnandB[23]), .ZN(AandB[23]) );
  NAND2_X1 U228 ( .A1(A[23]), .A2(B[23]), .ZN(AnandB[23]) );
  INV_X1 U229 ( .A(AnandB[22]), .ZN(AandB[22]) );
  NAND2_X1 U230 ( .A1(A[22]), .A2(B[22]), .ZN(AnandB[22]) );
  INV_X1 U231 ( .A(AnandB[21]), .ZN(AandB[21]) );
  NAND2_X1 U232 ( .A1(A[21]), .A2(B[21]), .ZN(AnandB[21]) );
  INV_X1 U233 ( .A(AnandB[20]), .ZN(AandB[20]) );
  NAND2_X1 U234 ( .A1(A[20]), .A2(B[20]), .ZN(AnandB[20]) );
  INV_X1 U235 ( .A(AnandB[18]), .ZN(AandB[18]) );
  NAND2_X1 U236 ( .A1(A[18]), .A2(B[18]), .ZN(AnandB[18]) );
  INV_X1 U237 ( .A(AnandB[17]), .ZN(AandB[17]) );
  NAND2_X1 U238 ( .A1(A[17]), .A2(B[17]), .ZN(AnandB[17]) );
  INV_X1 U239 ( .A(AnandB[16]), .ZN(AandB[16]) );
  NAND2_X1 U240 ( .A1(A[16]), .A2(B[16]), .ZN(AnandB[16]) );
  INV_X1 U241 ( .A(AnandB[6]), .ZN(AandB[6]) );
  NAND2_X1 U242 ( .A1(A[6]), .A2(B[6]), .ZN(AnandB[6]) );
  INV_X1 U243 ( .A(AnandB[5]), .ZN(AandB[5]) );
  NAND2_X1 U244 ( .A1(A[5]), .A2(B[5]), .ZN(AnandB[5]) );
  INV_X1 U245 ( .A(AnandB[4]), .ZN(AandB[4]) );
  NAND2_X1 U246 ( .A1(A[4]), .A2(B[4]), .ZN(AnandB[4]) );
  INV_X1 U247 ( .A(AnandB[12]), .ZN(AandB[12]) );
  NAND2_X1 U248 ( .A1(A[12]), .A2(B[12]), .ZN(AnandB[12]) );
  INV_X1 U249 ( .A(AnandB[11]), .ZN(AandB[11]) );
  NAND2_X1 U250 ( .A1(A[11]), .A2(B[11]), .ZN(AnandB[11]) );
  INV_X1 U251 ( .A(AnandB[10]), .ZN(AandB[10]) );
  NAND2_X1 U252 ( .A1(A[10]), .A2(B[10]), .ZN(AnandB[10]) );
  INV_X1 U253 ( .A(AnandB[9]), .ZN(AandB[9]) );
  NAND2_X1 U254 ( .A1(A[9]), .A2(B[9]), .ZN(AnandB[9]) );
  INV_X1 U255 ( .A(AnandB[7]), .ZN(AandB[7]) );
  NAND2_X1 U256 ( .A1(A[7]), .A2(B[7]), .ZN(AnandB[7]) );
endmodule


module Comp_Nbit32 ( signA, signB, Diff, Carry, unsign, AgB, AeqB, AnoteqB, 
        AlB, AgeqB, AleqB );
  input [31:0] Diff;
  input signA, signB, Carry, unsign;
  output AgB, AeqB, AnoteqB, AlB, AgeqB, AleqB;
  wire   n4, n6, n9, n10, n11, n12, n13, n14, n15, n16, n74, n76, n77, n79,
         n80, n81, n82;
  tri   unsign;

  NOR2_X1 U1 ( .A1(unsign), .A2(n6), .ZN(n4) );
  XOR2_X1 U2 ( .A(n74), .B(n4), .Z(AleqB) );
  XNOR2_X1 U3 ( .A(n82), .B(n4), .ZN(AgB) );
  NAND2_X1 U4 ( .A1(n79), .A2(Carry), .ZN(n74) );
  OR2_X1 U5 ( .A1(Diff[4]), .A2(Diff[5]), .ZN(n76) );
  NOR3_X1 U6 ( .A1(Diff[31]), .A2(Diff[3]), .A3(n76), .ZN(n15) );
  XNOR2_X1 U7 ( .A(Carry), .B(n4), .ZN(AlB) );
  NOR4_X1 U8 ( .A1(Diff[9]), .A2(Diff[8]), .A3(Diff[7]), .A4(Diff[6]), .ZN(n16) );
  XNOR2_X1 U9 ( .A(signB), .B(signA), .ZN(n6) );
  INV_X1 U10 ( .A(AlB), .ZN(AgeqB) );
  AND2_X1 U11 ( .A1(n9), .A2(n11), .ZN(n77) );
  AND3_X1 U12 ( .A1(n12), .A2(n10), .A3(n77), .ZN(n81) );
  NOR4_X1 U13 ( .A1(Diff[12]), .A2(Diff[11]), .A3(Diff[10]), .A4(Diff[0]), 
        .ZN(n9) );
  NOR4_X1 U14 ( .A1(Diff[16]), .A2(Diff[15]), .A3(Diff[14]), .A4(Diff[13]), 
        .ZN(n10) );
  NOR4_X1 U15 ( .A1(Diff[1]), .A2(Diff[19]), .A3(Diff[18]), .A4(Diff[17]), 
        .ZN(n11) );
  CLKBUF_X1 U16 ( .A(n79), .Z(AnoteqB) );
  INV_X1 U17 ( .A(AnoteqB), .ZN(AeqB) );
  NAND2_X1 U18 ( .A1(n80), .A2(n81), .ZN(n79) );
  AND4_X1 U19 ( .A1(n13), .A2(n16), .A3(n15), .A4(n14), .ZN(n80) );
  NOR4_X1 U20 ( .A1(Diff[23]), .A2(Diff[22]), .A3(Diff[21]), .A4(Diff[20]), 
        .ZN(n12) );
  NAND2_X1 U21 ( .A1(n79), .A2(Carry), .ZN(n82) );
  NOR4_X1 U22 ( .A1(Diff[30]), .A2(Diff[2]), .A3(Diff[29]), .A4(Diff[28]), 
        .ZN(n14) );
  NOR4_X1 U23 ( .A1(Diff[27]), .A2(Diff[26]), .A3(Diff[25]), .A4(Diff[24]), 
        .ZN(n13) );
endmodule


module AddSubN_Nbit32_1 ( A, B, addnsub, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input addnsub;
  output Cout;
  wire   n36, n42, n43, n44, n73, n77, n79, n86, n88, n95, n96, n99, net291417,
         net299273, net299291, net299504, n108, n112, net347328, net347340,
         net347354, net347489, net347504, net347548, n127, n138, net396670,
         net396766, net397095, net397133, net398565, n154, n158, n165, n176,
         n177, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201;
  wire   [31:0] addendB;
  wire   [7:0] Carry;
  assign n77 = A[3];
  assign n108 = A[9];
  assign n112 = A[5];
  assign n127 = A[1];
  assign n154 = A[0];
  assign n158 = addnsub;
  assign n176 = A[13];
  assign n177 = A[15];

  SparseTreeCarryGenN_Nbit32_1 STCG ( .A({A[31:16], n177, A[14], n176, 
        A[12:10], n108, A[8:6], n112, A[4], n77, A[2], n127, n154}), .B({
        addendB[31:29], n73, n86, addendB[26], n42, n165, n99, net347504, 
        net347548, n88, net347354, n43, n79, n138, net396766, net299273, 
        net397095, n36, net299291, net299504, net397133, n95, net347340, n96, 
        net347328, n44, net347489, net396670, net398565, net291417}), .Cin(
        n200), .Cout({Cout, Carry}) );
  CarrySumN_Nbit32_1 CSN ( .A({A[31:16], n177, A[14], n176, A[12:10], n108, 
        A[8:6], n112, A[4], n77, A[2], n127, n154}), .B({addendB[31:29], n73, 
        n86, addendB[26], n42, n165, n186, net347504, n182, n88, net347354, 
        n43, n79, n138, net396766, net299273, n187, n36, n189, n184, n185, n95, 
        n183, n188, n196, n44, n192, n190, n191, n197}), .Ci(Carry), .S(S) );
  XOR2_X1 U5 ( .A(n199), .B(B[8]), .Z(n95) );
  XOR2_X1 U7 ( .A(n199), .B(B[28]), .Z(n73) );
  XOR2_X1 U14 ( .A(n199), .B(B[22]), .Z(net347504) );
  XOR2_X1 U17 ( .A(n199), .B(B[10]), .Z(net299504) );
  XOR2_X1 U22 ( .A(n199), .B(B[27]), .Z(n86) );
  XOR2_X1 U24 ( .A(n199), .B(B[12]), .Z(n36) );
  XOR2_X1 U26 ( .A(n201), .B(B[20]), .Z(n88) );
  XOR2_X1 U27 ( .A(n201), .B(B[16]), .Z(n138) );
  XOR2_X1 U28 ( .A(n201), .B(B[24]), .Z(n165) );
  XOR2_X1 U29 ( .A(n201), .B(B[31]), .Z(addendB[31]) );
  XOR2_X1 U30 ( .A(n201), .B(B[30]), .Z(addendB[30]) );
  XOR2_X1 U31 ( .A(n201), .B(B[29]), .Z(addendB[29]) );
  XOR2_X1 U32 ( .A(n201), .B(B[26]), .Z(addendB[26]) );
  CLKBUF_X1 U1 ( .A(net347548), .Z(n182) );
  CLKBUF_X1 U2 ( .A(net347340), .Z(n183) );
  XNOR2_X1 U3 ( .A(n198), .B(B[7]), .ZN(net347340) );
  CLKBUF_X1 U4 ( .A(net299504), .Z(n184) );
  BUF_X1 U6 ( .A(n200), .Z(n199) );
  CLKBUF_X1 U8 ( .A(net397133), .Z(n185) );
  CLKBUF_X1 U9 ( .A(n99), .Z(n186) );
  CLKBUF_X1 U10 ( .A(net397095), .Z(n187) );
  CLKBUF_X1 U11 ( .A(n96), .Z(n188) );
  CLKBUF_X1 U12 ( .A(net299291), .Z(n189) );
  CLKBUF_X1 U13 ( .A(net396670), .Z(n190) );
  XOR2_X1 U15 ( .A(n199), .B(B[2]), .Z(net396670) );
  XNOR2_X1 U16 ( .A(B[0]), .B(n198), .ZN(n197) );
  CLKBUF_X1 U18 ( .A(net398565), .Z(n191) );
  XNOR2_X1 U19 ( .A(n198), .B(B[1]), .ZN(net398565) );
  XOR2_X1 U20 ( .A(n199), .B(B[25]), .Z(n42) );
  XOR2_X1 U21 ( .A(n199), .B(B[18]), .Z(n43) );
  XOR2_X1 U23 ( .A(n199), .B(B[17]), .Z(n79) );
  XOR2_X1 U25 ( .A(n199), .B(B[23]), .Z(n99) );
  XOR2_X1 U33 ( .A(B[5]), .B(n199), .Z(net347328) );
  NAND2_X1 U34 ( .A1(n194), .A2(n195), .ZN(net299291) );
  XOR2_X1 U35 ( .A(n199), .B(B[4]), .Z(n44) );
  XOR2_X1 U36 ( .A(n199), .B(B[6]), .Z(n96) );
  XNOR2_X1 U37 ( .A(n198), .B(B[14]), .ZN(net299273) );
  INV_X1 U38 ( .A(n199), .ZN(n198) );
  XOR2_X1 U39 ( .A(n199), .B(B[9]), .Z(net397133) );
  XOR2_X1 U40 ( .A(n199), .B(B[21]), .Z(net347548) );
  XOR2_X1 U41 ( .A(n199), .B(B[15]), .Z(net396766) );
  BUF_X1 U42 ( .A(n158), .Z(n200) );
  BUF_X1 U43 ( .A(n158), .Z(n201) );
  XOR2_X1 U44 ( .A(n199), .B(B[13]), .Z(net397095) );
  CLKBUF_X1 U45 ( .A(net347489), .Z(n192) );
  XNOR2_X1 U46 ( .A(B[3]), .B(n198), .ZN(net347489) );
  NAND2_X1 U47 ( .A1(n198), .A2(B[11]), .ZN(n194) );
  NAND2_X1 U48 ( .A1(n158), .A2(n193), .ZN(n195) );
  INV_X1 U49 ( .A(B[11]), .ZN(n193) );
  XOR2_X1 U50 ( .A(n199), .B(B[19]), .Z(net347354) );
  CLKBUF_X1 U51 ( .A(net347328), .Z(n196) );
  XNOR2_X1 U52 ( .A(B[0]), .B(n198), .ZN(net291417) );
endmodule


module BoothMulWallace_Nbit32 ( a, b, p );
  input [15:0] a;
  input [15:0] b;
  output [31:0] p;
  wire   init_0_0_port, init_0_1_port, init_0_2_port, init_0_3_port,
         init_0_4_port, init_0_5_port, init_0_6_port, init_0_7_port,
         init_0_8_port, init_0_9_port, init_0_10_port, init_0_11_port,
         init_0_12_port, init_0_13_port, init_0_14_port, init_1_1_port,
         init_1_2_port, init_1_3_port, init_1_4_port, init_1_5_port,
         init_1_6_port, init_1_7_port, init_1_8_port, init_1_9_port,
         init_1_10_port, init_1_11_port, init_1_12_port, init_1_13_port,
         init_1_14_port, init_1_15_port, init_2_2_port, init_2_3_port,
         init_2_4_port, init_2_5_port, init_2_6_port, init_2_7_port,
         init_2_8_port, init_2_9_port, init_2_10_port, init_2_11_port,
         init_2_12_port, init_2_13_port, init_2_14_port, init_2_15_port,
         init_2_16_port, first_out_0_0_port, first_out_0_1_port,
         first_out_0_2_port, first_out_0_3_port, first_out_0_4_port,
         first_out_0_5_port, first_out_0_6_port, first_out_0_7_port,
         first_out_0_8_port, first_out_0_9_port, first_out_0_10_port,
         first_out_0_11_port, first_out_0_12_port, first_out_0_13_port,
         first_out_0_14_port, first_out_0_15_port, first_out_0_16_port,
         first_out_0_17_port, first_out_0_18_port, first_out_0_19_port,
         first_out_0_20_port, first_out_0_21_port, first_out_0_22_port,
         first_out_0_23_port, first_out_0_24_port, first_out_0_25_port,
         first_out_0_26_port, first_out_0_27_port, first_out_0_28_port,
         first_out_0_29_port, first_out_0_30_port, first_out_0_31_port,
         first_cout_0_1_port, first_cout_0_2_port, first_cout_0_3_port,
         first_cout_0_4_port, first_cout_0_5_port, first_cout_0_6_port,
         first_cout_0_7_port, first_cout_0_8_port, first_cout_0_9_port,
         first_cout_0_10_port, first_cout_0_11_port, first_cout_0_12_port,
         first_cout_0_13_port, first_cout_0_14_port, first_cout_0_15_port,
         first_cout_0_16_port, first_cout_0_17_port, first_cout_0_18_port,
         first_cout_0_19_port, first_cout_0_20_port, first_cout_0_21_port,
         first_cout_0_22_port, first_cout_0_23_port, first_cout_0_24_port,
         first_cout_0_25_port, first_cout_0_26_port, first_cout_0_27_port,
         first_cout_0_28_port, first_cout_0_29_port, first_cout_0_30_port,
         first_cout_0_31_port, init_3_3_port, init_3_4_port, init_3_5_port,
         init_3_6_port, init_3_7_port, init_3_8_port, init_3_9_port,
         init_3_10_port, init_3_11_port, init_3_12_port, init_3_13_port,
         init_3_14_port, init_3_15_port, init_3_16_port, init_3_17_port,
         init_4_4_port, init_4_5_port, init_4_6_port, init_4_7_port,
         init_4_8_port, init_4_9_port, init_4_10_port, init_4_11_port,
         init_4_12_port, init_4_13_port, init_4_14_port, init_4_15_port,
         init_4_16_port, init_4_17_port, init_4_18_port, n443, init_5_5_port,
         init_5_6_port, init_5_7_port, init_5_8_port, init_5_9_port,
         init_5_10_port, init_5_11_port, init_5_12_port, init_5_13_port,
         init_5_14_port, init_5_15_port, init_5_16_port, init_5_17_port,
         init_5_18_port, init_5_19_port, init_5_31_port, first_out_1_0_port,
         first_out_1_1_port, first_out_1_2_port, first_out_1_3_port,
         first_out_1_4_port, first_out_1_5_port, first_out_1_6_port,
         first_out_1_7_port, first_out_1_8_port, first_out_1_9_port,
         first_out_1_10_port, first_out_1_11_port, first_out_1_12_port,
         first_out_1_13_port, first_out_1_14_port, first_out_1_15_port,
         first_out_1_16_port, first_out_1_17_port, first_out_1_18_port,
         first_out_1_19_port, first_out_1_20_port, first_out_1_21_port,
         first_out_1_22_port, first_out_1_23_port, first_out_1_24_port,
         first_out_1_25_port, first_out_1_26_port, first_out_1_27_port,
         first_out_1_28_port, first_out_1_29_port, first_out_1_30_port,
         first_out_1_31_port, first_cout_1_1_port, first_cout_1_2_port,
         first_cout_1_3_port, first_cout_1_4_port, first_cout_1_5_port,
         first_cout_1_6_port, first_cout_1_7_port, first_cout_1_8_port,
         first_cout_1_9_port, first_cout_1_10_port, first_cout_1_11_port,
         first_cout_1_12_port, first_cout_1_13_port, first_cout_1_14_port,
         first_cout_1_15_port, first_cout_1_16_port, first_cout_1_17_port,
         first_cout_1_18_port, first_cout_1_19_port, first_cout_1_20_port,
         first_cout_1_21_port, first_cout_1_22_port, first_cout_1_23_port,
         first_cout_1_24_port, first_cout_1_25_port, first_cout_1_26_port,
         first_cout_1_27_port, first_cout_1_28_port, first_cout_1_29_port,
         first_cout_1_30_port, first_cout_1_31_port, init_6_6_port,
         init_6_7_port, init_6_8_port, init_6_9_port, init_6_10_port,
         init_6_11_port, init_6_12_port, init_6_13_port, init_6_14_port,
         init_6_15_port, init_6_16_port, init_6_17_port, init_6_18_port,
         init_6_19_port, init_6_20_port, n431, init_7_7_port, init_7_8_port,
         init_7_9_port, init_7_10_port, init_7_11_port, init_7_12_port,
         init_7_13_port, init_7_14_port, init_7_15_port, init_7_16_port,
         init_7_17_port, init_7_18_port, init_7_19_port, init_7_20_port,
         init_7_21_port, n425, init_8_8_port, init_8_9_port, init_8_10_port,
         init_8_11_port, init_8_12_port, init_8_13_port, init_8_14_port,
         init_8_15_port, init_8_16_port, init_8_17_port, init_8_18_port,
         init_8_19_port, init_8_20_port, init_8_21_port, init_8_22_port,
         init_8_31_port, first_out_2_0_port, first_out_2_1_port,
         first_out_2_2_port, first_out_2_3_port, first_out_2_4_port,
         first_out_2_5_port, first_out_2_6_port, first_out_2_7_port,
         first_out_2_8_port, first_out_2_9_port, first_out_2_10_port,
         first_out_2_11_port, first_out_2_12_port, first_out_2_13_port,
         first_out_2_14_port, first_out_2_15_port, first_out_2_16_port,
         first_out_2_17_port, first_out_2_18_port, first_out_2_19_port,
         first_out_2_20_port, first_out_2_21_port, first_out_2_22_port,
         first_out_2_23_port, first_out_2_24_port, first_out_2_25_port,
         first_out_2_26_port, first_out_2_27_port, first_out_2_28_port,
         first_out_2_29_port, first_out_2_30_port, first_out_2_31_port,
         first_cout_2_1_port, first_cout_2_2_port, first_cout_2_3_port,
         first_cout_2_4_port, first_cout_2_5_port, first_cout_2_6_port,
         first_cout_2_7_port, first_cout_2_8_port, first_cout_2_9_port,
         first_cout_2_10_port, first_cout_2_11_port, first_cout_2_12_port,
         first_cout_2_13_port, first_cout_2_14_port, first_cout_2_15_port,
         first_cout_2_16_port, first_cout_2_17_port, first_cout_2_18_port,
         first_cout_2_19_port, first_cout_2_20_port, first_cout_2_21_port,
         first_cout_2_22_port, first_cout_2_23_port, first_cout_2_24_port,
         first_cout_2_25_port, first_cout_2_26_port, first_cout_2_27_port,
         first_cout_2_28_port, first_cout_2_29_port, first_cout_2_30_port,
         first_cout_2_31_port, init_9_9_port, init_9_10_port, init_9_11_port,
         init_9_12_port, init_9_13_port, init_9_14_port, init_9_15_port,
         init_9_16_port, init_9_17_port, init_9_18_port, init_9_19_port,
         init_9_20_port, init_9_21_port, init_9_22_port, init_9_23_port, n418,
         init_10_10_port, init_10_11_port, init_10_12_port, init_10_13_port,
         init_10_14_port, init_10_15_port, init_10_16_port, init_10_17_port,
         init_10_18_port, init_10_19_port, init_10_20_port, init_10_21_port,
         init_10_22_port, init_10_23_port, init_10_24_port, n420,
         init_11_11_port, init_11_12_port, init_11_13_port, init_11_14_port,
         init_11_15_port, init_11_16_port, init_11_17_port, init_11_18_port,
         init_11_19_port, init_11_20_port, init_11_21_port, init_11_22_port,
         init_11_23_port, init_11_24_port, init_11_25_port, n411,
         first_out_3_0_port, first_out_3_1_port, first_out_3_2_port,
         first_out_3_3_port, first_out_3_4_port, first_out_3_5_port,
         first_out_3_6_port, first_out_3_7_port, first_out_3_8_port,
         first_out_3_9_port, first_out_3_10_port, first_out_3_11_port,
         first_out_3_12_port, first_out_3_13_port, first_out_3_14_port,
         first_out_3_15_port, first_out_3_16_port, first_out_3_17_port,
         first_out_3_18_port, first_out_3_19_port, first_out_3_20_port,
         first_out_3_21_port, first_out_3_22_port, first_out_3_23_port,
         first_out_3_24_port, first_out_3_25_port, first_out_3_26_port,
         first_out_3_27_port, first_out_3_28_port, first_out_3_29_port,
         first_out_3_30_port, first_out_3_31_port, first_cout_3_1_port,
         first_cout_3_2_port, first_cout_3_3_port, first_cout_3_4_port,
         first_cout_3_5_port, first_cout_3_6_port, first_cout_3_7_port,
         first_cout_3_8_port, first_cout_3_9_port, first_cout_3_10_port,
         first_cout_3_11_port, first_cout_3_12_port, first_cout_3_13_port,
         first_cout_3_14_port, first_cout_3_15_port, first_cout_3_16_port,
         first_cout_3_17_port, first_cout_3_18_port, first_cout_3_19_port,
         first_cout_3_20_port, first_cout_3_21_port, first_cout_3_22_port,
         first_cout_3_23_port, first_cout_3_24_port, first_cout_3_25_port,
         first_cout_3_26_port, first_cout_3_27_port, first_cout_3_28_port,
         first_cout_3_29_port, first_cout_3_30_port, first_cout_3_31_port,
         init_12_12_port, init_12_13_port, init_12_14_port, init_12_15_port,
         init_12_16_port, init_12_17_port, init_12_18_port, init_12_19_port,
         init_12_20_port, init_12_21_port, init_12_22_port, init_12_23_port,
         init_12_24_port, init_12_25_port, init_12_26_port, init_12_31_port,
         init_13_13_port, init_13_14_port, init_13_15_port, init_13_16_port,
         init_13_17_port, init_13_18_port, init_13_19_port, init_13_20_port,
         init_13_21_port, init_13_22_port, init_13_23_port, init_13_24_port,
         init_13_25_port, init_13_26_port, init_13_27_port, init_13_31_port,
         init_14_14_port, init_14_15_port, init_14_16_port, init_14_17_port,
         init_14_18_port, init_14_19_port, init_14_20_port, init_14_21_port,
         init_14_22_port, init_14_23_port, init_14_24_port, init_14_25_port,
         init_14_26_port, init_14_27_port, init_14_28_port, init_14_31_port,
         first_out_4_0_port, first_out_4_1_port, first_out_4_2_port,
         first_out_4_3_port, first_out_4_4_port, first_out_4_5_port,
         first_out_4_6_port, first_out_4_7_port, first_out_4_8_port,
         first_out_4_9_port, first_out_4_10_port, first_out_4_11_port,
         first_out_4_12_port, first_out_4_13_port, first_out_4_14_port,
         first_out_4_15_port, first_out_4_16_port, first_out_4_17_port,
         first_out_4_18_port, first_out_4_19_port, first_out_4_20_port,
         first_out_4_21_port, first_out_4_22_port, first_out_4_23_port,
         first_out_4_24_port, first_out_4_25_port, first_out_4_26_port,
         first_out_4_27_port, first_out_4_28_port, first_out_4_29_port,
         first_out_4_30_port, first_out_4_31_port, first_cout_4_1_port,
         first_cout_4_2_port, first_cout_4_3_port, first_cout_4_4_port,
         first_cout_4_5_port, first_cout_4_6_port, first_cout_4_7_port,
         first_cout_4_8_port, first_cout_4_9_port, first_cout_4_10_port,
         first_cout_4_11_port, first_cout_4_12_port, first_cout_4_13_port,
         first_cout_4_14_port, first_cout_4_15_port, first_cout_4_16_port,
         first_cout_4_17_port, first_cout_4_18_port, first_cout_4_19_port,
         first_cout_4_20_port, first_cout_4_21_port, first_cout_4_22_port,
         first_cout_4_23_port, first_cout_4_24_port, first_cout_4_25_port,
         first_cout_4_26_port, first_cout_4_27_port, first_cout_4_28_port,
         first_cout_4_29_port, first_cout_4_30_port, first_cout_4_31_port,
         second_out_0_0_port, second_out_0_1_port, second_out_0_2_port,
         second_out_0_3_port, second_out_0_4_port, second_out_0_5_port,
         second_out_0_6_port, second_out_0_7_port, second_out_0_8_port,
         second_out_0_9_port, second_out_0_10_port, second_out_0_11_port,
         second_out_0_12_port, second_out_0_13_port, second_out_0_14_port,
         second_out_0_15_port, second_out_0_16_port, second_out_0_17_port,
         second_out_0_18_port, second_out_0_19_port, second_out_0_20_port,
         second_out_0_21_port, second_out_0_22_port, second_out_0_23_port,
         second_out_0_24_port, second_out_0_25_port, second_out_0_26_port,
         second_out_0_27_port, second_out_0_28_port, second_out_0_29_port,
         second_out_0_30_port, second_out_0_31_port, second_cout_0_1_port,
         second_cout_0_2_port, second_cout_0_3_port, second_cout_0_4_port,
         second_cout_0_5_port, second_cout_0_6_port, second_cout_0_7_port,
         second_cout_0_8_port, second_cout_0_9_port, second_cout_0_10_port,
         second_cout_0_11_port, second_cout_0_12_port, second_cout_0_13_port,
         second_cout_0_14_port, second_cout_0_15_port, second_cout_0_16_port,
         second_cout_0_17_port, second_cout_0_18_port, second_cout_0_19_port,
         second_cout_0_20_port, second_cout_0_21_port, second_cout_0_22_port,
         second_cout_0_23_port, second_cout_0_24_port, second_cout_0_25_port,
         second_cout_0_26_port, second_cout_0_27_port, second_cout_0_28_port,
         second_cout_0_29_port, second_cout_0_30_port, second_cout_0_31_port,
         second_out_1_0_port, second_out_1_1_port, second_out_1_2_port,
         second_out_1_3_port, second_out_1_4_port, second_out_1_5_port,
         second_out_1_6_port, second_out_1_7_port, second_out_1_8_port,
         second_out_1_9_port, second_out_1_10_port, second_out_1_11_port,
         second_out_1_12_port, second_out_1_13_port, second_out_1_14_port,
         second_out_1_15_port, second_out_1_16_port, second_out_1_17_port,
         second_out_1_18_port, second_out_1_19_port, second_out_1_20_port,
         second_out_1_21_port, second_out_1_22_port, second_out_1_23_port,
         second_out_1_24_port, second_out_1_25_port, second_out_1_26_port,
         second_out_1_27_port, second_out_1_28_port, second_out_1_29_port,
         second_out_1_30_port, second_out_1_31_port, second_cout_1_1_port,
         second_cout_1_2_port, second_cout_1_3_port, second_cout_1_4_port,
         second_cout_1_5_port, second_cout_1_6_port, second_cout_1_7_port,
         second_cout_1_8_port, second_cout_1_9_port, second_cout_1_10_port,
         second_cout_1_11_port, second_cout_1_12_port, second_cout_1_13_port,
         second_cout_1_14_port, second_cout_1_15_port, second_cout_1_16_port,
         second_cout_1_17_port, second_cout_1_18_port, second_cout_1_19_port,
         second_cout_1_20_port, second_cout_1_21_port, second_cout_1_22_port,
         second_cout_1_23_port, second_cout_1_24_port, second_cout_1_25_port,
         second_cout_1_26_port, second_cout_1_27_port, second_cout_1_28_port,
         second_cout_1_29_port, second_cout_1_30_port, second_cout_1_31_port,
         second_out_2_0_port, second_out_2_1_port, second_out_2_2_port,
         second_out_2_3_port, second_out_2_4_port, second_out_2_5_port,
         second_out_2_6_port, second_out_2_7_port, second_out_2_8_port,
         second_out_2_9_port, second_out_2_10_port, second_out_2_11_port,
         second_out_2_12_port, second_out_2_13_port, second_out_2_14_port,
         second_out_2_15_port, second_out_2_16_port, second_out_2_17_port,
         second_out_2_18_port, second_out_2_19_port, second_out_2_20_port,
         second_out_2_21_port, second_out_2_22_port, second_out_2_23_port,
         second_out_2_24_port, second_out_2_25_port, second_out_2_26_port,
         second_out_2_27_port, second_out_2_28_port, second_out_2_29_port,
         second_out_2_30_port, second_out_2_31_port, second_cout_2_1_port,
         second_cout_2_2_port, second_cout_2_3_port, second_cout_2_4_port,
         second_cout_2_5_port, second_cout_2_6_port, second_cout_2_7_port,
         second_cout_2_8_port, second_cout_2_9_port, second_cout_2_10_port,
         second_cout_2_11_port, second_cout_2_12_port, second_cout_2_13_port,
         second_cout_2_14_port, second_cout_2_15_port, second_cout_2_16_port,
         second_cout_2_17_port, second_cout_2_18_port, second_cout_2_19_port,
         second_cout_2_20_port, second_cout_2_21_port, second_cout_2_22_port,
         second_cout_2_23_port, second_cout_2_24_port, second_cout_2_25_port,
         second_cout_2_26_port, second_cout_2_27_port, second_cout_2_28_port,
         second_cout_2_29_port, second_cout_2_30_port, second_cout_2_31_port,
         third_out_0_0_port, third_out_0_1_port, third_out_0_2_port,
         third_out_0_3_port, third_out_0_4_port, third_out_0_5_port,
         third_out_0_6_port, third_out_0_7_port, third_out_0_8_port,
         third_out_0_9_port, third_out_0_10_port, third_out_0_11_port,
         third_out_0_12_port, third_out_0_13_port, third_out_0_14_port,
         third_out_0_15_port, third_out_0_16_port, third_out_0_17_port,
         third_out_0_18_port, third_out_0_19_port, third_out_0_20_port,
         third_out_0_21_port, third_out_0_22_port, third_out_0_23_port,
         third_out_0_24_port, third_out_0_25_port, third_out_0_26_port,
         third_out_0_27_port, third_out_0_28_port, third_out_0_29_port,
         third_out_0_30_port, third_out_0_31_port, third_cout_0_1_port,
         third_cout_0_2_port, third_cout_0_3_port, third_cout_0_4_port,
         third_cout_0_5_port, third_cout_0_6_port, third_cout_0_7_port,
         third_cout_0_8_port, third_cout_0_9_port, third_cout_0_10_port,
         third_cout_0_11_port, third_cout_0_12_port, third_cout_0_13_port,
         third_cout_0_14_port, third_cout_0_15_port, third_cout_0_16_port,
         third_cout_0_17_port, third_cout_0_18_port, third_cout_0_19_port,
         third_cout_0_20_port, third_cout_0_21_port, third_cout_0_22_port,
         third_cout_0_23_port, third_cout_0_24_port, third_cout_0_25_port,
         third_cout_0_26_port, third_cout_0_27_port, third_cout_0_28_port,
         third_cout_0_29_port, third_cout_0_30_port, third_cout_0_31_port,
         third_out_1_0_port, third_out_1_1_port, third_out_1_2_port,
         third_out_1_3_port, third_out_1_4_port, third_out_1_5_port,
         third_out_1_6_port, third_out_1_7_port, third_out_1_8_port,
         third_out_1_9_port, third_out_1_10_port, third_out_1_11_port,
         third_out_1_12_port, third_out_1_13_port, third_out_1_14_port,
         third_out_1_15_port, third_out_1_16_port, third_out_1_17_port,
         third_out_1_18_port, third_out_1_19_port, third_out_1_20_port,
         third_out_1_21_port, third_out_1_22_port, third_out_1_23_port,
         third_out_1_24_port, third_out_1_25_port, third_out_1_26_port,
         third_out_1_27_port, third_out_1_28_port, third_out_1_29_port,
         third_out_1_30_port, third_out_1_31_port, third_cout_1_1_port,
         third_cout_1_2_port, third_cout_1_3_port, third_cout_1_4_port,
         third_cout_1_5_port, third_cout_1_6_port, third_cout_1_7_port,
         third_cout_1_8_port, third_cout_1_9_port, third_cout_1_10_port,
         third_cout_1_11_port, third_cout_1_12_port, third_cout_1_13_port,
         third_cout_1_14_port, third_cout_1_15_port, third_cout_1_16_port,
         third_cout_1_17_port, third_cout_1_18_port, third_cout_1_19_port,
         third_cout_1_20_port, third_cout_1_21_port, third_cout_1_22_port,
         third_cout_1_23_port, third_cout_1_24_port, third_cout_1_25_port,
         third_cout_1_26_port, third_cout_1_27_port, third_cout_1_28_port,
         third_cout_1_29_port, third_cout_1_30_port, third_cout_1_31_port,
         fourth_out_0_0_port, fourth_out_0_1_port, fourth_out_0_2_port,
         fourth_out_0_3_port, fourth_out_0_4_port, fourth_out_0_5_port,
         fourth_out_0_6_port, fourth_out_0_7_port, fourth_out_0_8_port,
         fourth_out_0_9_port, fourth_out_0_10_port, fourth_out_0_11_port,
         fourth_out_0_12_port, fourth_out_0_13_port, fourth_out_0_14_port,
         fourth_out_0_15_port, fourth_out_0_16_port, fourth_out_0_17_port,
         fourth_out_0_18_port, fourth_out_0_19_port, fourth_out_0_20_port,
         fourth_out_0_21_port, fourth_out_0_22_port, fourth_out_0_23_port,
         fourth_out_0_24_port, fourth_out_0_25_port, fourth_out_0_26_port,
         fourth_out_0_27_port, fourth_out_0_28_port, fourth_out_0_29_port,
         fourth_out_0_30_port, fourth_out_0_31_port, fourth_cout_0_1_port,
         fourth_cout_0_2_port, fourth_cout_0_3_port, fourth_cout_0_4_port,
         fourth_cout_0_5_port, fourth_cout_0_6_port, fourth_cout_0_7_port,
         fourth_cout_0_8_port, fourth_cout_0_9_port, fourth_cout_0_10_port,
         fourth_cout_0_11_port, fourth_cout_0_12_port, fourth_cout_0_13_port,
         fourth_cout_0_14_port, fourth_cout_0_15_port, fourth_cout_0_16_port,
         fourth_cout_0_17_port, fourth_cout_0_18_port, fourth_cout_0_19_port,
         fourth_cout_0_20_port, fourth_cout_0_21_port, fourth_cout_0_22_port,
         fourth_cout_0_23_port, fourth_cout_0_24_port, fourth_cout_0_25_port,
         fourth_cout_0_26_port, fourth_cout_0_27_port, fourth_cout_0_28_port,
         fourth_cout_0_29_port, fourth_cout_0_30_port, fourth_cout_0_31_port,
         init_15_15_port, init_15_16_port, init_15_17_port, init_15_18_port,
         init_15_19_port, init_15_20_port, n409, n410, init_15_23_port,
         init_15_24_port, init_15_25_port, init_15_26_port, init_15_27_port,
         init_15_28_port, init_15_29_port, init_15_31_port,
         fourth_out_1_0_port, fourth_out_1_1_port, fourth_out_1_2_port,
         fourth_out_1_3_port, fourth_out_1_4_port, fourth_out_1_5_port,
         fourth_out_1_6_port, fourth_out_1_7_port, fourth_out_1_8_port,
         fourth_out_1_9_port, fourth_out_1_10_port, fourth_out_1_11_port,
         fourth_out_1_12_port, fourth_out_1_13_port, fourth_out_1_14_port,
         fourth_out_1_15_port, fourth_out_1_16_port, fourth_out_1_17_port,
         fourth_out_1_18_port, fourth_out_1_19_port, fourth_out_1_20_port,
         fourth_out_1_21_port, fourth_out_1_22_port, fourth_out_1_23_port,
         fourth_out_1_24_port, fourth_out_1_25_port, fourth_out_1_26_port,
         fourth_out_1_27_port, fourth_out_1_28_port, fourth_out_1_29_port,
         fourth_out_1_30_port, fourth_out_1_31_port, fourth_cout_1_1_port,
         fourth_cout_1_2_port, fourth_cout_1_3_port, fourth_cout_1_4_port,
         fourth_cout_1_5_port, fourth_cout_1_6_port, fourth_cout_1_7_port,
         fourth_cout_1_8_port, fourth_cout_1_9_port, fourth_cout_1_10_port,
         fourth_cout_1_11_port, fourth_cout_1_12_port, fourth_cout_1_13_port,
         fourth_cout_1_14_port, fourth_cout_1_15_port, fourth_cout_1_16_port,
         fourth_cout_1_17_port, fourth_cout_1_18_port, fourth_cout_1_19_port,
         fourth_cout_1_20_port, fourth_cout_1_21_port, fourth_cout_1_22_port,
         fourth_cout_1_23_port, fourth_cout_1_24_port, fourth_cout_1_25_port,
         fourth_cout_1_26_port, fourth_cout_1_27_port, fourth_cout_1_28_port,
         fourth_cout_1_29_port, fourth_cout_1_30_port, fourth_cout_1_31_port,
         fifth_out_0_port, fifth_out_1_port, fifth_out_2_port,
         fifth_out_3_port, fifth_out_4_port, fifth_out_5_port,
         fifth_out_6_port, fifth_out_7_port, fifth_out_8_port,
         fifth_out_9_port, fifth_out_10_port, fifth_out_11_port,
         fifth_out_12_port, fifth_out_13_port, fifth_out_14_port,
         fifth_out_15_port, fifth_out_16_port, fifth_out_17_port,
         fifth_out_18_port, fifth_out_19_port, fifth_out_20_port,
         fifth_out_21_port, fifth_out_22_port, fifth_out_23_port,
         fifth_out_24_port, fifth_out_25_port, fifth_out_26_port,
         fifth_out_27_port, fifth_out_28_port, fifth_out_29_port,
         fifth_out_30_port, fifth_out_31_port, fifth_cout_1_port,
         fifth_cout_2_port, fifth_cout_3_port, fifth_cout_4_port,
         fifth_cout_5_port, fifth_cout_6_port, fifth_cout_7_port,
         fifth_cout_8_port, fifth_cout_9_port, fifth_cout_10_port,
         fifth_cout_11_port, fifth_cout_12_port, fifth_cout_13_port,
         fifth_cout_14_port, fifth_cout_15_port, fifth_cout_16_port,
         fifth_cout_17_port, fifth_cout_18_port, fifth_cout_19_port,
         fifth_cout_20_port, fifth_cout_21_port, fifth_cout_22_port,
         fifth_cout_23_port, fifth_cout_24_port, fifth_cout_25_port,
         fifth_cout_26_port, fifth_cout_27_port, fifth_cout_28_port,
         fifth_cout_29_port, fifth_cout_30_port, fifth_cout_31_port,
         sixth_out_0_port, sixth_out_1_port, sixth_out_2_port,
         sixth_out_3_port, sixth_out_4_port, sixth_out_5_port,
         sixth_out_6_port, sixth_out_7_port, sixth_out_8_port,
         sixth_out_9_port, sixth_out_10_port, sixth_out_11_port,
         sixth_out_12_port, sixth_out_13_port, sixth_out_14_port,
         sixth_out_15_port, sixth_out_16_port, sixth_out_17_port,
         sixth_out_18_port, sixth_out_19_port, sixth_out_20_port,
         sixth_out_21_port, sixth_out_22_port, sixth_out_23_port,
         sixth_out_24_port, sixth_out_25_port, sixth_out_26_port,
         sixth_out_27_port, sixth_out_28_port, sixth_out_29_port,
         sixth_out_30_port, sixth_out_31_port, sixth_cout_1_port,
         sixth_cout_2_port, sixth_cout_3_port, sixth_cout_4_port,
         sixth_cout_5_port, sixth_cout_6_port, sixth_cout_7_port,
         sixth_cout_8_port, sixth_cout_9_port, sixth_cout_10_port,
         sixth_cout_11_port, sixth_cout_12_port, sixth_cout_13_port,
         sixth_cout_14_port, sixth_cout_15_port, sixth_cout_16_port,
         sixth_cout_17_port, sixth_cout_18_port, sixth_cout_19_port,
         sixth_cout_20_port, sixth_cout_21_port, sixth_cout_22_port,
         sixth_cout_23_port, sixth_cout_24_port, sixth_cout_25_port,
         sixth_cout_26_port, sixth_cout_27_port, sixth_cout_28_port,
         sixth_cout_29_port, sixth_cout_30_port, sixth_cout_31_port, N49, N48,
         N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N132,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, n247, n248, n249, n250, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n102, n103, n104, n105, n106, n107, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13;

  CSA_N32_0 CSA0 ( .A({n258, n258, n258, n258, n258, n257, n257, n257, n257, 
        n257, n257, n257, n257, n257, n257, n257, n257, init_0_14_port, 
        init_0_13_port, init_0_12_port, init_0_11_port, init_0_10_port, 
        init_0_9_port, init_0_8_port, init_0_7_port, init_0_6_port, 
        init_0_5_port, init_0_4_port, init_0_3_port, init_0_2_port, 
        init_0_1_port, init_0_0_port}), .B({n260, n260, n260, n260, n259, n259, 
        n259, n259, n259, n259, n259, n259, n259, n259, n259, n259, 
        init_1_15_port, init_1_14_port, init_1_13_port, init_1_12_port, 
        init_1_11_port, init_1_10_port, init_1_9_port, init_1_8_port, 
        init_1_7_port, init_1_6_port, init_1_5_port, init_1_4_port, 
        init_1_3_port, init_1_2_port, init_1_1_port, 1'b0}), .C({n262, n262, 
        n262, n261, n261, n261, n261, n261, n261, n261, n261, n261, n261, n261, 
        n261, init_2_16_port, init_2_15_port, init_2_14_port, init_2_13_port, 
        init_2_12_port, init_2_11_port, init_2_10_port, init_2_9_port, 
        init_2_8_port, init_2_7_port, init_2_6_port, init_2_5_port, 
        init_2_4_port, init_2_3_port, init_2_2_port, 1'b0, 1'b0}), .sum_out({
        first_out_0_31_port, first_out_0_30_port, first_out_0_29_port, 
        first_out_0_28_port, first_out_0_27_port, first_out_0_26_port, 
        first_out_0_25_port, first_out_0_24_port, first_out_0_23_port, 
        first_out_0_22_port, first_out_0_21_port, first_out_0_20_port, 
        first_out_0_19_port, first_out_0_18_port, first_out_0_17_port, 
        first_out_0_16_port, first_out_0_15_port, first_out_0_14_port, 
        first_out_0_13_port, first_out_0_12_port, first_out_0_11_port, 
        first_out_0_10_port, first_out_0_9_port, first_out_0_8_port, 
        first_out_0_7_port, first_out_0_6_port, first_out_0_5_port, 
        first_out_0_4_port, first_out_0_3_port, first_out_0_2_port, 
        first_out_0_1_port, first_out_0_0_port}), .cout({first_cout_0_31_port, 
        first_cout_0_30_port, first_cout_0_29_port, first_cout_0_28_port, 
        first_cout_0_27_port, first_cout_0_26_port, first_cout_0_25_port, 
        first_cout_0_24_port, first_cout_0_23_port, first_cout_0_22_port, 
        first_cout_0_21_port, first_cout_0_20_port, first_cout_0_19_port, 
        first_cout_0_18_port, first_cout_0_17_port, first_cout_0_16_port, 
        first_cout_0_15_port, first_cout_0_14_port, first_cout_0_13_port, 
        first_cout_0_12_port, first_cout_0_11_port, first_cout_0_10_port, 
        first_cout_0_9_port, first_cout_0_8_port, first_cout_0_7_port, 
        first_cout_0_6_port, first_cout_0_5_port, first_cout_0_4_port, 
        first_cout_0_3_port, first_cout_0_2_port, first_cout_0_1_port, 
        SYNOPSYS_UNCONNECTED__0}) );
  CSA_N32_13 CSA1 ( .A({n264, n264, n263, n263, n263, n263, n263, n263, n263, 
        n263, n263, n263, n263, n263, init_3_17_port, init_3_16_port, 
        init_3_15_port, init_3_14_port, init_3_13_port, init_3_12_port, 
        init_3_11_port, init_3_10_port, init_3_9_port, init_3_8_port, 
        init_3_7_port, init_3_6_port, init_3_5_port, init_3_4_port, 
        init_3_3_port, 1'b0, 1'b0, 1'b0}), .B({n443, n266, n266, n266, n266, 
        n266, n266, n265, n265, n265, n265, n265, n265, init_4_18_port, 
        init_4_17_port, init_4_16_port, init_4_15_port, init_4_14_port, 
        init_4_13_port, init_4_12_port, init_4_11_port, init_4_10_port, 
        init_4_9_port, init_4_8_port, init_4_7_port, init_4_6_port, 
        init_4_5_port, init_4_4_port, 1'b0, 1'b0, 1'b0, 1'b0}), .C({
        init_5_31_port, init_5_31_port, init_5_31_port, init_5_31_port, 
        init_5_31_port, init_5_31_port, init_5_31_port, init_5_31_port, 
        init_5_31_port, init_5_31_port, init_5_31_port, init_5_31_port, 
        init_5_19_port, init_5_18_port, init_5_17_port, init_5_16_port, 
        init_5_15_port, init_5_14_port, init_5_13_port, init_5_12_port, 
        init_5_11_port, init_5_10_port, init_5_9_port, init_5_8_port, 
        init_5_7_port, init_5_6_port, init_5_5_port, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .sum_out({first_out_1_31_port, first_out_1_30_port, 
        first_out_1_29_port, first_out_1_28_port, first_out_1_27_port, 
        first_out_1_26_port, first_out_1_25_port, first_out_1_24_port, 
        first_out_1_23_port, first_out_1_22_port, first_out_1_21_port, 
        first_out_1_20_port, first_out_1_19_port, first_out_1_18_port, 
        first_out_1_17_port, first_out_1_16_port, first_out_1_15_port, 
        first_out_1_14_port, first_out_1_13_port, first_out_1_12_port, 
        first_out_1_11_port, first_out_1_10_port, first_out_1_9_port, 
        first_out_1_8_port, first_out_1_7_port, first_out_1_6_port, 
        first_out_1_5_port, first_out_1_4_port, first_out_1_3_port, 
        first_out_1_2_port, first_out_1_1_port, first_out_1_0_port}), .cout({
        first_cout_1_31_port, first_cout_1_30_port, first_cout_1_29_port, 
        first_cout_1_28_port, first_cout_1_27_port, first_cout_1_26_port, 
        first_cout_1_25_port, first_cout_1_24_port, first_cout_1_23_port, 
        first_cout_1_22_port, first_cout_1_21_port, first_cout_1_20_port, 
        first_cout_1_19_port, first_cout_1_18_port, first_cout_1_17_port, 
        first_cout_1_16_port, first_cout_1_15_port, first_cout_1_14_port, 
        first_cout_1_13_port, first_cout_1_12_port, first_cout_1_11_port, 
        first_cout_1_10_port, first_cout_1_9_port, first_cout_1_8_port, 
        first_cout_1_7_port, first_cout_1_6_port, first_cout_1_5_port, 
        first_cout_1_4_port, first_cout_1_3_port, first_cout_1_2_port, 
        first_cout_1_1_port, SYNOPSYS_UNCONNECTED__1}) );
  CSA_N32_12 CSA2 ( .A({n431, n431, n431, n431, n431, n431, n431, n431, n431, 
        n431, n431, init_6_20_port, init_6_19_port, init_6_18_port, 
        init_6_17_port, init_6_16_port, init_6_15_port, init_6_14_port, 
        init_6_13_port, init_6_12_port, init_6_11_port, init_6_10_port, 
        init_6_9_port, init_6_8_port, init_6_7_port, init_6_6_port, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({n425, n425, n425, n425, n425, n425, n425, 
        n425, n425, n425, init_7_21_port, init_7_20_port, init_7_19_port, 
        init_7_18_port, init_7_17_port, init_7_16_port, init_7_15_port, 
        init_7_14_port, init_7_13_port, init_7_12_port, init_7_11_port, 
        init_7_10_port, init_7_9_port, init_7_8_port, init_7_7_port, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({init_8_31_port, 
        init_8_31_port, init_8_31_port, init_8_31_port, init_8_31_port, 
        init_8_31_port, init_8_31_port, init_8_31_port, init_8_31_port, 
        init_8_22_port, init_8_21_port, init_8_20_port, init_8_19_port, 
        init_8_18_port, init_8_17_port, init_8_16_port, init_8_15_port, 
        init_8_14_port, init_8_13_port, init_8_12_port, init_8_11_port, 
        init_8_10_port, init_8_9_port, init_8_8_port, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .sum_out({first_out_2_31_port, 
        first_out_2_30_port, first_out_2_29_port, first_out_2_28_port, 
        first_out_2_27_port, first_out_2_26_port, first_out_2_25_port, 
        first_out_2_24_port, first_out_2_23_port, first_out_2_22_port, 
        first_out_2_21_port, first_out_2_20_port, first_out_2_19_port, 
        first_out_2_18_port, first_out_2_17_port, first_out_2_16_port, 
        first_out_2_15_port, first_out_2_14_port, first_out_2_13_port, 
        first_out_2_12_port, first_out_2_11_port, first_out_2_10_port, 
        first_out_2_9_port, first_out_2_8_port, first_out_2_7_port, 
        first_out_2_6_port, first_out_2_5_port, first_out_2_4_port, 
        first_out_2_3_port, first_out_2_2_port, first_out_2_1_port, 
        first_out_2_0_port}), .cout({first_cout_2_31_port, 
        first_cout_2_30_port, first_cout_2_29_port, first_cout_2_28_port, 
        first_cout_2_27_port, first_cout_2_26_port, first_cout_2_25_port, 
        first_cout_2_24_port, first_cout_2_23_port, first_cout_2_22_port, 
        first_cout_2_21_port, first_cout_2_20_port, first_cout_2_19_port, 
        first_cout_2_18_port, first_cout_2_17_port, first_cout_2_16_port, 
        first_cout_2_15_port, first_cout_2_14_port, first_cout_2_13_port, 
        first_cout_2_12_port, first_cout_2_11_port, first_cout_2_10_port, 
        first_cout_2_9_port, first_cout_2_8_port, first_cout_2_7_port, 
        first_cout_2_6_port, first_cout_2_5_port, first_cout_2_4_port, 
        first_cout_2_3_port, first_cout_2_2_port, first_cout_2_1_port, 
        SYNOPSYS_UNCONNECTED__2}) );
  CSA_N32_11 CSA3 ( .A({n418, n418, n418, n418, n418, n418, n418, n418, 
        init_9_23_port, init_9_22_port, init_9_21_port, init_9_20_port, 
        init_9_19_port, init_9_18_port, init_9_17_port, init_9_16_port, 
        init_9_15_port, init_9_14_port, init_9_13_port, init_9_12_port, 
        init_9_11_port, init_9_10_port, init_9_9_port, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n420, n420, n420, n420, n420, n420, 
        n420, init_10_24_port, init_10_23_port, init_10_22_port, 
        init_10_21_port, init_10_20_port, init_10_19_port, init_10_18_port, 
        init_10_17_port, init_10_16_port, init_10_15_port, init_10_14_port, 
        init_10_13_port, init_10_12_port, init_10_11_port, init_10_10_port, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({n411, 
        n411, n411, n411, n411, n411, init_11_25_port, init_11_24_port, 
        init_11_23_port, init_11_22_port, init_11_21_port, init_11_20_port, 
        init_11_19_port, init_11_18_port, init_11_17_port, init_11_16_port, 
        init_11_15_port, init_11_14_port, init_11_13_port, init_11_12_port, 
        init_11_11_port, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .sum_out({first_out_3_31_port, first_out_3_30_port, 
        first_out_3_29_port, first_out_3_28_port, first_out_3_27_port, 
        first_out_3_26_port, first_out_3_25_port, first_out_3_24_port, 
        first_out_3_23_port, first_out_3_22_port, first_out_3_21_port, 
        first_out_3_20_port, first_out_3_19_port, first_out_3_18_port, 
        first_out_3_17_port, first_out_3_16_port, first_out_3_15_port, 
        first_out_3_14_port, first_out_3_13_port, first_out_3_12_port, 
        first_out_3_11_port, first_out_3_10_port, first_out_3_9_port, 
        first_out_3_8_port, first_out_3_7_port, first_out_3_6_port, 
        first_out_3_5_port, first_out_3_4_port, first_out_3_3_port, 
        first_out_3_2_port, first_out_3_1_port, first_out_3_0_port}), .cout({
        first_cout_3_31_port, first_cout_3_30_port, first_cout_3_29_port, 
        first_cout_3_28_port, first_cout_3_27_port, first_cout_3_26_port, 
        first_cout_3_25_port, first_cout_3_24_port, first_cout_3_23_port, 
        first_cout_3_22_port, first_cout_3_21_port, first_cout_3_20_port, 
        first_cout_3_19_port, first_cout_3_18_port, first_cout_3_17_port, 
        first_cout_3_16_port, first_cout_3_15_port, first_cout_3_14_port, 
        first_cout_3_13_port, first_cout_3_12_port, first_cout_3_11_port, 
        first_cout_3_10_port, first_cout_3_9_port, first_cout_3_8_port, 
        first_cout_3_7_port, first_cout_3_6_port, first_cout_3_5_port, 
        first_cout_3_4_port, first_cout_3_3_port, first_cout_3_2_port, 
        first_cout_3_1_port, SYNOPSYS_UNCONNECTED__3}) );
  CSA_N32_10 CSA4 ( .A({init_12_31_port, init_12_31_port, init_12_31_port, 
        init_12_31_port, init_12_31_port, init_12_26_port, init_12_25_port, 
        init_12_24_port, init_12_23_port, init_12_22_port, init_12_21_port, 
        init_12_20_port, init_12_19_port, init_12_18_port, init_12_17_port, 
        init_12_16_port, init_12_15_port, init_12_14_port, init_12_13_port, 
        init_12_12_port, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({init_13_31_port, init_13_31_port, 
        init_13_31_port, init_13_31_port, init_13_27_port, init_13_26_port, 
        init_13_25_port, init_13_24_port, init_13_23_port, init_13_22_port, 
        init_13_21_port, init_13_20_port, init_13_19_port, init_13_18_port, 
        init_13_17_port, init_13_16_port, init_13_15_port, init_13_14_port, 
        init_13_13_port, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .C({init_14_31_port, init_14_31_port, 
        init_14_31_port, init_14_28_port, init_14_27_port, init_14_26_port, 
        init_14_25_port, init_14_24_port, init_14_23_port, init_14_22_port, 
        init_14_21_port, init_14_20_port, init_14_19_port, init_14_18_port, 
        init_14_17_port, init_14_16_port, init_14_15_port, init_14_14_port, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .sum_out({first_out_4_31_port, first_out_4_30_port, 
        first_out_4_29_port, first_out_4_28_port, first_out_4_27_port, 
        first_out_4_26_port, first_out_4_25_port, first_out_4_24_port, 
        first_out_4_23_port, first_out_4_22_port, first_out_4_21_port, 
        first_out_4_20_port, first_out_4_19_port, first_out_4_18_port, 
        first_out_4_17_port, first_out_4_16_port, first_out_4_15_port, 
        first_out_4_14_port, first_out_4_13_port, first_out_4_12_port, 
        first_out_4_11_port, first_out_4_10_port, first_out_4_9_port, 
        first_out_4_8_port, first_out_4_7_port, first_out_4_6_port, 
        first_out_4_5_port, first_out_4_4_port, first_out_4_3_port, 
        first_out_4_2_port, first_out_4_1_port, first_out_4_0_port}), .cout({
        first_cout_4_31_port, first_cout_4_30_port, first_cout_4_29_port, 
        first_cout_4_28_port, first_cout_4_27_port, first_cout_4_26_port, 
        first_cout_4_25_port, first_cout_4_24_port, first_cout_4_23_port, 
        first_cout_4_22_port, first_cout_4_21_port, first_cout_4_20_port, 
        first_cout_4_19_port, first_cout_4_18_port, first_cout_4_17_port, 
        first_cout_4_16_port, first_cout_4_15_port, first_cout_4_14_port, 
        first_cout_4_13_port, first_cout_4_12_port, first_cout_4_11_port, 
        first_cout_4_10_port, first_cout_4_9_port, first_cout_4_8_port, 
        first_cout_4_7_port, first_cout_4_6_port, first_cout_4_5_port, 
        first_cout_4_4_port, first_cout_4_3_port, first_cout_4_2_port, 
        first_cout_4_1_port, SYNOPSYS_UNCONNECTED__4}) );
  CSA_N32_9 CSA5 ( .A({first_out_0_31_port, first_out_0_30_port, 
        first_out_0_29_port, first_out_0_28_port, first_out_0_27_port, 
        first_out_0_26_port, first_out_0_25_port, first_out_0_24_port, 
        first_out_0_23_port, first_out_0_22_port, first_out_0_21_port, 
        first_out_0_20_port, first_out_0_19_port, first_out_0_18_port, 
        first_out_0_17_port, first_out_0_16_port, first_out_0_15_port, 
        first_out_0_14_port, first_out_0_13_port, first_out_0_12_port, 
        first_out_0_11_port, first_out_0_10_port, first_out_0_9_port, 
        first_out_0_8_port, first_out_0_7_port, first_out_0_6_port, 
        first_out_0_5_port, first_out_0_4_port, first_out_0_3_port, 
        first_out_0_2_port, first_out_0_1_port, first_out_0_0_port}), .B({
        first_cout_0_31_port, first_cout_0_30_port, first_cout_0_29_port, 
        first_cout_0_28_port, first_cout_0_27_port, first_cout_0_26_port, 
        first_cout_0_25_port, first_cout_0_24_port, first_cout_0_23_port, 
        first_cout_0_22_port, first_cout_0_21_port, first_cout_0_20_port, 
        first_cout_0_19_port, first_cout_0_18_port, first_cout_0_17_port, 
        first_cout_0_16_port, first_cout_0_15_port, first_cout_0_14_port, 
        first_cout_0_13_port, first_cout_0_12_port, first_cout_0_11_port, 
        first_cout_0_10_port, first_cout_0_9_port, first_cout_0_8_port, 
        first_cout_0_7_port, first_cout_0_6_port, first_cout_0_5_port, 
        first_cout_0_4_port, first_cout_0_3_port, first_cout_0_2_port, 
        first_cout_0_1_port, 1'b0}), .C({first_out_1_31_port, 
        first_out_1_30_port, first_out_1_29_port, first_out_1_28_port, 
        first_out_1_27_port, first_out_1_26_port, first_out_1_25_port, 
        first_out_1_24_port, first_out_1_23_port, first_out_1_22_port, 
        first_out_1_21_port, first_out_1_20_port, first_out_1_19_port, 
        first_out_1_18_port, first_out_1_17_port, first_out_1_16_port, 
        first_out_1_15_port, first_out_1_14_port, first_out_1_13_port, 
        first_out_1_12_port, first_out_1_11_port, first_out_1_10_port, 
        first_out_1_9_port, first_out_1_8_port, first_out_1_7_port, 
        first_out_1_6_port, first_out_1_5_port, first_out_1_4_port, 
        first_out_1_3_port, first_out_1_2_port, first_out_1_1_port, 
        first_out_1_0_port}), .sum_out({second_out_0_31_port, 
        second_out_0_30_port, second_out_0_29_port, second_out_0_28_port, 
        second_out_0_27_port, second_out_0_26_port, second_out_0_25_port, 
        second_out_0_24_port, second_out_0_23_port, second_out_0_22_port, 
        second_out_0_21_port, second_out_0_20_port, second_out_0_19_port, 
        second_out_0_18_port, second_out_0_17_port, second_out_0_16_port, 
        second_out_0_15_port, second_out_0_14_port, second_out_0_13_port, 
        second_out_0_12_port, second_out_0_11_port, second_out_0_10_port, 
        second_out_0_9_port, second_out_0_8_port, second_out_0_7_port, 
        second_out_0_6_port, second_out_0_5_port, second_out_0_4_port, 
        second_out_0_3_port, second_out_0_2_port, second_out_0_1_port, 
        second_out_0_0_port}), .cout({second_cout_0_31_port, 
        second_cout_0_30_port, second_cout_0_29_port, second_cout_0_28_port, 
        second_cout_0_27_port, second_cout_0_26_port, second_cout_0_25_port, 
        second_cout_0_24_port, second_cout_0_23_port, second_cout_0_22_port, 
        second_cout_0_21_port, second_cout_0_20_port, second_cout_0_19_port, 
        second_cout_0_18_port, second_cout_0_17_port, second_cout_0_16_port, 
        second_cout_0_15_port, second_cout_0_14_port, second_cout_0_13_port, 
        second_cout_0_12_port, second_cout_0_11_port, second_cout_0_10_port, 
        second_cout_0_9_port, second_cout_0_8_port, second_cout_0_7_port, 
        second_cout_0_6_port, second_cout_0_5_port, second_cout_0_4_port, 
        second_cout_0_3_port, second_cout_0_2_port, second_cout_0_1_port, 
        SYNOPSYS_UNCONNECTED__5}) );
  CSA_N32_8 CSA6 ( .A({first_cout_1_31_port, first_cout_1_30_port, 
        first_cout_1_29_port, first_cout_1_28_port, first_cout_1_27_port, 
        first_cout_1_26_port, first_cout_1_25_port, first_cout_1_24_port, 
        first_cout_1_23_port, first_cout_1_22_port, first_cout_1_21_port, 
        first_cout_1_20_port, first_cout_1_19_port, first_cout_1_18_port, 
        first_cout_1_17_port, first_cout_1_16_port, first_cout_1_15_port, 
        first_cout_1_14_port, first_cout_1_13_port, first_cout_1_12_port, 
        first_cout_1_11_port, first_cout_1_10_port, first_cout_1_9_port, 
        first_cout_1_8_port, first_cout_1_7_port, first_cout_1_6_port, 
        first_cout_1_5_port, first_cout_1_4_port, first_cout_1_3_port, 
        first_cout_1_2_port, first_cout_1_1_port, 1'b0}), .B({
        first_out_2_31_port, first_out_2_30_port, first_out_2_29_port, 
        first_out_2_28_port, first_out_2_27_port, first_out_2_26_port, 
        first_out_2_25_port, first_out_2_24_port, first_out_2_23_port, 
        first_out_2_22_port, first_out_2_21_port, first_out_2_20_port, 
        first_out_2_19_port, first_out_2_18_port, first_out_2_17_port, 
        first_out_2_16_port, first_out_2_15_port, first_out_2_14_port, 
        first_out_2_13_port, first_out_2_12_port, first_out_2_11_port, 
        first_out_2_10_port, first_out_2_9_port, first_out_2_8_port, 
        first_out_2_7_port, first_out_2_6_port, first_out_2_5_port, 
        first_out_2_4_port, first_out_2_3_port, first_out_2_2_port, 
        first_out_2_1_port, first_out_2_0_port}), .C({first_cout_2_31_port, 
        first_cout_2_30_port, first_cout_2_29_port, first_cout_2_28_port, 
        first_cout_2_27_port, first_cout_2_26_port, first_cout_2_25_port, 
        first_cout_2_24_port, first_cout_2_23_port, first_cout_2_22_port, 
        first_cout_2_21_port, first_cout_2_20_port, first_cout_2_19_port, 
        first_cout_2_18_port, first_cout_2_17_port, first_cout_2_16_port, 
        first_cout_2_15_port, first_cout_2_14_port, first_cout_2_13_port, 
        first_cout_2_12_port, first_cout_2_11_port, first_cout_2_10_port, 
        first_cout_2_9_port, first_cout_2_8_port, first_cout_2_7_port, 
        first_cout_2_6_port, first_cout_2_5_port, first_cout_2_4_port, 
        first_cout_2_3_port, first_cout_2_2_port, first_cout_2_1_port, 1'b0}), 
        .sum_out({second_out_1_31_port, second_out_1_30_port, 
        second_out_1_29_port, second_out_1_28_port, second_out_1_27_port, 
        second_out_1_26_port, second_out_1_25_port, second_out_1_24_port, 
        second_out_1_23_port, second_out_1_22_port, second_out_1_21_port, 
        second_out_1_20_port, second_out_1_19_port, second_out_1_18_port, 
        second_out_1_17_port, second_out_1_16_port, second_out_1_15_port, 
        second_out_1_14_port, second_out_1_13_port, second_out_1_12_port, 
        second_out_1_11_port, second_out_1_10_port, second_out_1_9_port, 
        second_out_1_8_port, second_out_1_7_port, second_out_1_6_port, 
        second_out_1_5_port, second_out_1_4_port, second_out_1_3_port, 
        second_out_1_2_port, second_out_1_1_port, second_out_1_0_port}), 
        .cout({second_cout_1_31_port, second_cout_1_30_port, 
        second_cout_1_29_port, second_cout_1_28_port, second_cout_1_27_port, 
        second_cout_1_26_port, second_cout_1_25_port, second_cout_1_24_port, 
        second_cout_1_23_port, second_cout_1_22_port, second_cout_1_21_port, 
        second_cout_1_20_port, second_cout_1_19_port, second_cout_1_18_port, 
        second_cout_1_17_port, second_cout_1_16_port, second_cout_1_15_port, 
        second_cout_1_14_port, second_cout_1_13_port, second_cout_1_12_port, 
        second_cout_1_11_port, second_cout_1_10_port, second_cout_1_9_port, 
        second_cout_1_8_port, second_cout_1_7_port, second_cout_1_6_port, 
        second_cout_1_5_port, second_cout_1_4_port, second_cout_1_3_port, 
        second_cout_1_2_port, second_cout_1_1_port, SYNOPSYS_UNCONNECTED__6})
         );
  CSA_N32_7 CSA7 ( .A({first_out_3_31_port, first_out_3_30_port, 
        first_out_3_29_port, first_out_3_28_port, first_out_3_27_port, 
        first_out_3_26_port, first_out_3_25_port, first_out_3_24_port, 
        first_out_3_23_port, first_out_3_22_port, first_out_3_21_port, 
        first_out_3_20_port, first_out_3_19_port, first_out_3_18_port, 
        first_out_3_17_port, first_out_3_16_port, first_out_3_15_port, 
        first_out_3_14_port, first_out_3_13_port, first_out_3_12_port, 
        first_out_3_11_port, first_out_3_10_port, first_out_3_9_port, 
        first_out_3_8_port, first_out_3_7_port, first_out_3_6_port, 
        first_out_3_5_port, first_out_3_4_port, first_out_3_3_port, 
        first_out_3_2_port, first_out_3_1_port, first_out_3_0_port}), .B({
        first_cout_3_31_port, first_cout_3_30_port, first_cout_3_29_port, 
        first_cout_3_28_port, first_cout_3_27_port, first_cout_3_26_port, 
        first_cout_3_25_port, first_cout_3_24_port, first_cout_3_23_port, 
        first_cout_3_22_port, first_cout_3_21_port, first_cout_3_20_port, 
        first_cout_3_19_port, first_cout_3_18_port, first_cout_3_17_port, 
        first_cout_3_16_port, first_cout_3_15_port, first_cout_3_14_port, 
        first_cout_3_13_port, first_cout_3_12_port, first_cout_3_11_port, 
        first_cout_3_10_port, first_cout_3_9_port, first_cout_3_8_port, 
        first_cout_3_7_port, first_cout_3_6_port, first_cout_3_5_port, 
        first_cout_3_4_port, first_cout_3_3_port, first_cout_3_2_port, 
        first_cout_3_1_port, 1'b0}), .C({first_out_4_31_port, 
        first_out_4_30_port, first_out_4_29_port, first_out_4_28_port, 
        first_out_4_27_port, first_out_4_26_port, first_out_4_25_port, 
        first_out_4_24_port, first_out_4_23_port, first_out_4_22_port, 
        first_out_4_21_port, first_out_4_20_port, first_out_4_19_port, 
        first_out_4_18_port, first_out_4_17_port, first_out_4_16_port, 
        first_out_4_15_port, first_out_4_14_port, first_out_4_13_port, 
        first_out_4_12_port, first_out_4_11_port, first_out_4_10_port, 
        first_out_4_9_port, first_out_4_8_port, first_out_4_7_port, 
        first_out_4_6_port, first_out_4_5_port, first_out_4_4_port, 
        first_out_4_3_port, first_out_4_2_port, first_out_4_1_port, 
        first_out_4_0_port}), .sum_out({second_out_2_31_port, 
        second_out_2_30_port, second_out_2_29_port, second_out_2_28_port, 
        second_out_2_27_port, second_out_2_26_port, second_out_2_25_port, 
        second_out_2_24_port, second_out_2_23_port, second_out_2_22_port, 
        second_out_2_21_port, second_out_2_20_port, second_out_2_19_port, 
        second_out_2_18_port, second_out_2_17_port, second_out_2_16_port, 
        second_out_2_15_port, second_out_2_14_port, second_out_2_13_port, 
        second_out_2_12_port, second_out_2_11_port, second_out_2_10_port, 
        second_out_2_9_port, second_out_2_8_port, second_out_2_7_port, 
        second_out_2_6_port, second_out_2_5_port, second_out_2_4_port, 
        second_out_2_3_port, second_out_2_2_port, second_out_2_1_port, 
        second_out_2_0_port}), .cout({second_cout_2_31_port, 
        second_cout_2_30_port, second_cout_2_29_port, second_cout_2_28_port, 
        second_cout_2_27_port, second_cout_2_26_port, second_cout_2_25_port, 
        second_cout_2_24_port, second_cout_2_23_port, second_cout_2_22_port, 
        second_cout_2_21_port, second_cout_2_20_port, second_cout_2_19_port, 
        second_cout_2_18_port, second_cout_2_17_port, second_cout_2_16_port, 
        second_cout_2_15_port, second_cout_2_14_port, second_cout_2_13_port, 
        second_cout_2_12_port, second_cout_2_11_port, second_cout_2_10_port, 
        second_cout_2_9_port, second_cout_2_8_port, second_cout_2_7_port, 
        second_cout_2_6_port, second_cout_2_5_port, second_cout_2_4_port, 
        second_cout_2_3_port, second_cout_2_2_port, second_cout_2_1_port, 
        SYNOPSYS_UNCONNECTED__7}) );
  CSA_N32_6 CSA8 ( .A({second_out_0_31_port, second_out_0_30_port, 
        second_out_0_29_port, second_out_0_28_port, second_out_0_27_port, 
        second_out_0_26_port, second_out_0_25_port, second_out_0_24_port, 
        second_out_0_23_port, second_out_0_22_port, second_out_0_21_port, 
        second_out_0_20_port, second_out_0_19_port, second_out_0_18_port, 
        second_out_0_17_port, second_out_0_16_port, second_out_0_15_port, 
        second_out_0_14_port, second_out_0_13_port, second_out_0_12_port, 
        second_out_0_11_port, second_out_0_10_port, second_out_0_9_port, 
        second_out_0_8_port, second_out_0_7_port, second_out_0_6_port, 
        second_out_0_5_port, second_out_0_4_port, second_out_0_3_port, 
        second_out_0_2_port, second_out_0_1_port, second_out_0_0_port}), .B({
        second_cout_0_31_port, second_cout_0_30_port, second_cout_0_29_port, 
        second_cout_0_28_port, second_cout_0_27_port, second_cout_0_26_port, 
        second_cout_0_25_port, second_cout_0_24_port, second_cout_0_23_port, 
        second_cout_0_22_port, second_cout_0_21_port, second_cout_0_20_port, 
        second_cout_0_19_port, second_cout_0_18_port, second_cout_0_17_port, 
        second_cout_0_16_port, second_cout_0_15_port, second_cout_0_14_port, 
        second_cout_0_13_port, second_cout_0_12_port, second_cout_0_11_port, 
        second_cout_0_10_port, second_cout_0_9_port, second_cout_0_8_port, 
        second_cout_0_7_port, second_cout_0_6_port, second_cout_0_5_port, 
        second_cout_0_4_port, second_cout_0_3_port, second_cout_0_2_port, 
        second_cout_0_1_port, 1'b0}), .C({second_out_1_31_port, 
        second_out_1_30_port, second_out_1_29_port, second_out_1_28_port, 
        second_out_1_27_port, second_out_1_26_port, second_out_1_25_port, 
        second_out_1_24_port, second_out_1_23_port, second_out_1_22_port, 
        second_out_1_21_port, second_out_1_20_port, second_out_1_19_port, 
        second_out_1_18_port, second_out_1_17_port, second_out_1_16_port, 
        second_out_1_15_port, second_out_1_14_port, second_out_1_13_port, 
        second_out_1_12_port, second_out_1_11_port, second_out_1_10_port, 
        second_out_1_9_port, second_out_1_8_port, second_out_1_7_port, 
        second_out_1_6_port, second_out_1_5_port, second_out_1_4_port, 
        second_out_1_3_port, second_out_1_2_port, second_out_1_1_port, 
        second_out_1_0_port}), .sum_out({third_out_0_31_port, 
        third_out_0_30_port, third_out_0_29_port, third_out_0_28_port, 
        third_out_0_27_port, third_out_0_26_port, third_out_0_25_port, 
        third_out_0_24_port, third_out_0_23_port, third_out_0_22_port, 
        third_out_0_21_port, third_out_0_20_port, third_out_0_19_port, 
        third_out_0_18_port, third_out_0_17_port, third_out_0_16_port, 
        third_out_0_15_port, third_out_0_14_port, third_out_0_13_port, 
        third_out_0_12_port, third_out_0_11_port, third_out_0_10_port, 
        third_out_0_9_port, third_out_0_8_port, third_out_0_7_port, 
        third_out_0_6_port, third_out_0_5_port, third_out_0_4_port, 
        third_out_0_3_port, third_out_0_2_port, third_out_0_1_port, 
        third_out_0_0_port}), .cout({third_cout_0_31_port, 
        third_cout_0_30_port, third_cout_0_29_port, third_cout_0_28_port, 
        third_cout_0_27_port, third_cout_0_26_port, third_cout_0_25_port, 
        third_cout_0_24_port, third_cout_0_23_port, third_cout_0_22_port, 
        third_cout_0_21_port, third_cout_0_20_port, third_cout_0_19_port, 
        third_cout_0_18_port, third_cout_0_17_port, third_cout_0_16_port, 
        third_cout_0_15_port, third_cout_0_14_port, third_cout_0_13_port, 
        third_cout_0_12_port, third_cout_0_11_port, third_cout_0_10_port, 
        third_cout_0_9_port, third_cout_0_8_port, third_cout_0_7_port, 
        third_cout_0_6_port, third_cout_0_5_port, third_cout_0_4_port, 
        third_cout_0_3_port, third_cout_0_2_port, third_cout_0_1_port, 
        SYNOPSYS_UNCONNECTED__8}) );
  CSA_N32_5 CSA9 ( .A({second_cout_1_31_port, second_cout_1_30_port, 
        second_cout_1_29_port, second_cout_1_28_port, second_cout_1_27_port, 
        second_cout_1_26_port, second_cout_1_25_port, second_cout_1_24_port, 
        second_cout_1_23_port, second_cout_1_22_port, second_cout_1_21_port, 
        second_cout_1_20_port, second_cout_1_19_port, second_cout_1_18_port, 
        second_cout_1_17_port, second_cout_1_16_port, second_cout_1_15_port, 
        second_cout_1_14_port, second_cout_1_13_port, second_cout_1_12_port, 
        second_cout_1_11_port, second_cout_1_10_port, second_cout_1_9_port, 
        second_cout_1_8_port, second_cout_1_7_port, second_cout_1_6_port, 
        second_cout_1_5_port, second_cout_1_4_port, second_cout_1_3_port, 
        second_cout_1_2_port, second_cout_1_1_port, 1'b0}), .B({
        second_out_2_31_port, second_out_2_30_port, second_out_2_29_port, 
        second_out_2_28_port, second_out_2_27_port, second_out_2_26_port, 
        second_out_2_25_port, second_out_2_24_port, second_out_2_23_port, 
        second_out_2_22_port, second_out_2_21_port, second_out_2_20_port, 
        second_out_2_19_port, second_out_2_18_port, second_out_2_17_port, 
        second_out_2_16_port, second_out_2_15_port, second_out_2_14_port, 
        second_out_2_13_port, second_out_2_12_port, second_out_2_11_port, 
        second_out_2_10_port, second_out_2_9_port, second_out_2_8_port, 
        second_out_2_7_port, second_out_2_6_port, second_out_2_5_port, 
        second_out_2_4_port, second_out_2_3_port, second_out_2_2_port, 
        second_out_2_1_port, second_out_2_0_port}), .C({second_cout_2_31_port, 
        second_cout_2_30_port, second_cout_2_29_port, second_cout_2_28_port, 
        second_cout_2_27_port, second_cout_2_26_port, second_cout_2_25_port, 
        second_cout_2_24_port, second_cout_2_23_port, second_cout_2_22_port, 
        second_cout_2_21_port, second_cout_2_20_port, second_cout_2_19_port, 
        second_cout_2_18_port, second_cout_2_17_port, second_cout_2_16_port, 
        second_cout_2_15_port, second_cout_2_14_port, second_cout_2_13_port, 
        second_cout_2_12_port, second_cout_2_11_port, second_cout_2_10_port, 
        second_cout_2_9_port, second_cout_2_8_port, second_cout_2_7_port, 
        second_cout_2_6_port, second_cout_2_5_port, second_cout_2_4_port, 
        second_cout_2_3_port, second_cout_2_2_port, second_cout_2_1_port, 1'b0}), .sum_out({third_out_1_31_port, third_out_1_30_port, third_out_1_29_port, 
        third_out_1_28_port, third_out_1_27_port, third_out_1_26_port, 
        third_out_1_25_port, third_out_1_24_port, third_out_1_23_port, 
        third_out_1_22_port, third_out_1_21_port, third_out_1_20_port, 
        third_out_1_19_port, third_out_1_18_port, third_out_1_17_port, 
        third_out_1_16_port, third_out_1_15_port, third_out_1_14_port, 
        third_out_1_13_port, third_out_1_12_port, third_out_1_11_port, 
        third_out_1_10_port, third_out_1_9_port, third_out_1_8_port, 
        third_out_1_7_port, third_out_1_6_port, third_out_1_5_port, 
        third_out_1_4_port, third_out_1_3_port, third_out_1_2_port, 
        third_out_1_1_port, third_out_1_0_port}), .cout({third_cout_1_31_port, 
        third_cout_1_30_port, third_cout_1_29_port, third_cout_1_28_port, 
        third_cout_1_27_port, third_cout_1_26_port, third_cout_1_25_port, 
        third_cout_1_24_port, third_cout_1_23_port, third_cout_1_22_port, 
        third_cout_1_21_port, third_cout_1_20_port, third_cout_1_19_port, 
        third_cout_1_18_port, third_cout_1_17_port, third_cout_1_16_port, 
        third_cout_1_15_port, third_cout_1_14_port, third_cout_1_13_port, 
        third_cout_1_12_port, third_cout_1_11_port, third_cout_1_10_port, 
        third_cout_1_9_port, third_cout_1_8_port, third_cout_1_7_port, 
        third_cout_1_6_port, third_cout_1_5_port, third_cout_1_4_port, 
        third_cout_1_3_port, third_cout_1_2_port, third_cout_1_1_port, 
        SYNOPSYS_UNCONNECTED__9}) );
  CSA_N32_4 CSA10 ( .A({third_out_0_31_port, third_out_0_30_port, 
        third_out_0_29_port, third_out_0_28_port, third_out_0_27_port, 
        third_out_0_26_port, third_out_0_25_port, third_out_0_24_port, 
        third_out_0_23_port, third_out_0_22_port, third_out_0_21_port, 
        third_out_0_20_port, third_out_0_19_port, third_out_0_18_port, 
        third_out_0_17_port, third_out_0_16_port, third_out_0_15_port, 
        third_out_0_14_port, third_out_0_13_port, third_out_0_12_port, 
        third_out_0_11_port, third_out_0_10_port, third_out_0_9_port, 
        third_out_0_8_port, third_out_0_7_port, third_out_0_6_port, 
        third_out_0_5_port, third_out_0_4_port, third_out_0_3_port, 
        third_out_0_2_port, third_out_0_1_port, third_out_0_0_port}), .B({
        third_cout_0_31_port, third_cout_0_30_port, third_cout_0_29_port, 
        third_cout_0_28_port, third_cout_0_27_port, third_cout_0_26_port, 
        third_cout_0_25_port, third_cout_0_24_port, third_cout_0_23_port, 
        third_cout_0_22_port, third_cout_0_21_port, third_cout_0_20_port, 
        third_cout_0_19_port, third_cout_0_18_port, third_cout_0_17_port, 
        third_cout_0_16_port, third_cout_0_15_port, third_cout_0_14_port, 
        third_cout_0_13_port, third_cout_0_12_port, third_cout_0_11_port, 
        third_cout_0_10_port, third_cout_0_9_port, third_cout_0_8_port, 
        third_cout_0_7_port, third_cout_0_6_port, third_cout_0_5_port, 
        third_cout_0_4_port, third_cout_0_3_port, third_cout_0_2_port, 
        third_cout_0_1_port, 1'b0}), .C({third_out_1_31_port, 
        third_out_1_30_port, third_out_1_29_port, third_out_1_28_port, 
        third_out_1_27_port, third_out_1_26_port, third_out_1_25_port, 
        third_out_1_24_port, third_out_1_23_port, third_out_1_22_port, 
        third_out_1_21_port, third_out_1_20_port, third_out_1_19_port, 
        third_out_1_18_port, third_out_1_17_port, third_out_1_16_port, 
        third_out_1_15_port, third_out_1_14_port, third_out_1_13_port, 
        third_out_1_12_port, third_out_1_11_port, third_out_1_10_port, 
        third_out_1_9_port, third_out_1_8_port, third_out_1_7_port, 
        third_out_1_6_port, third_out_1_5_port, third_out_1_4_port, 
        third_out_1_3_port, third_out_1_2_port, third_out_1_1_port, 
        third_out_1_0_port}), .sum_out({fourth_out_0_31_port, 
        fourth_out_0_30_port, fourth_out_0_29_port, fourth_out_0_28_port, 
        fourth_out_0_27_port, fourth_out_0_26_port, fourth_out_0_25_port, 
        fourth_out_0_24_port, fourth_out_0_23_port, fourth_out_0_22_port, 
        fourth_out_0_21_port, fourth_out_0_20_port, fourth_out_0_19_port, 
        fourth_out_0_18_port, fourth_out_0_17_port, fourth_out_0_16_port, 
        fourth_out_0_15_port, fourth_out_0_14_port, fourth_out_0_13_port, 
        fourth_out_0_12_port, fourth_out_0_11_port, fourth_out_0_10_port, 
        fourth_out_0_9_port, fourth_out_0_8_port, fourth_out_0_7_port, 
        fourth_out_0_6_port, fourth_out_0_5_port, fourth_out_0_4_port, 
        fourth_out_0_3_port, fourth_out_0_2_port, fourth_out_0_1_port, 
        fourth_out_0_0_port}), .cout({fourth_cout_0_31_port, 
        fourth_cout_0_30_port, fourth_cout_0_29_port, fourth_cout_0_28_port, 
        fourth_cout_0_27_port, fourth_cout_0_26_port, fourth_cout_0_25_port, 
        fourth_cout_0_24_port, fourth_cout_0_23_port, fourth_cout_0_22_port, 
        fourth_cout_0_21_port, fourth_cout_0_20_port, fourth_cout_0_19_port, 
        fourth_cout_0_18_port, fourth_cout_0_17_port, fourth_cout_0_16_port, 
        fourth_cout_0_15_port, fourth_cout_0_14_port, fourth_cout_0_13_port, 
        fourth_cout_0_12_port, fourth_cout_0_11_port, fourth_cout_0_10_port, 
        fourth_cout_0_9_port, fourth_cout_0_8_port, fourth_cout_0_7_port, 
        fourth_cout_0_6_port, fourth_cout_0_5_port, fourth_cout_0_4_port, 
        fourth_cout_0_3_port, fourth_cout_0_2_port, fourth_cout_0_1_port, 
        SYNOPSYS_UNCONNECTED__10}) );
  CSA_N32_3 CSA11 ( .A({third_cout_1_31_port, third_cout_1_30_port, 
        third_cout_1_29_port, third_cout_1_28_port, third_cout_1_27_port, 
        third_cout_1_26_port, third_cout_1_25_port, third_cout_1_24_port, 
        third_cout_1_23_port, third_cout_1_22_port, third_cout_1_21_port, 
        third_cout_1_20_port, third_cout_1_19_port, third_cout_1_18_port, 
        third_cout_1_17_port, third_cout_1_16_port, third_cout_1_15_port, 
        third_cout_1_14_port, third_cout_1_13_port, third_cout_1_12_port, 
        third_cout_1_11_port, third_cout_1_10_port, third_cout_1_9_port, 
        third_cout_1_8_port, third_cout_1_7_port, third_cout_1_6_port, 
        third_cout_1_5_port, third_cout_1_4_port, third_cout_1_3_port, 
        third_cout_1_2_port, third_cout_1_1_port, 1'b0}), .B({
        first_cout_4_31_port, first_cout_4_30_port, first_cout_4_29_port, 
        first_cout_4_28_port, first_cout_4_27_port, first_cout_4_26_port, 
        first_cout_4_25_port, first_cout_4_24_port, first_cout_4_23_port, 
        first_cout_4_22_port, first_cout_4_21_port, first_cout_4_20_port, 
        first_cout_4_19_port, first_cout_4_18_port, first_cout_4_17_port, 
        first_cout_4_16_port, first_cout_4_15_port, first_cout_4_14_port, 
        first_cout_4_13_port, first_cout_4_12_port, first_cout_4_11_port, 
        first_cout_4_10_port, first_cout_4_9_port, first_cout_4_8_port, 
        first_cout_4_7_port, first_cout_4_6_port, first_cout_4_5_port, 
        first_cout_4_4_port, first_cout_4_3_port, first_cout_4_2_port, 
        first_cout_4_1_port, 1'b0}), .C({init_15_31_port, init_15_31_port, 
        init_15_29_port, init_15_28_port, init_15_27_port, init_15_26_port, 
        init_15_25_port, init_15_24_port, init_15_23_port, n410, n409, 
        init_15_20_port, init_15_19_port, init_15_18_port, init_15_17_port, 
        init_15_16_port, init_15_15_port, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum_out({
        fourth_out_1_31_port, fourth_out_1_30_port, fourth_out_1_29_port, 
        fourth_out_1_28_port, fourth_out_1_27_port, fourth_out_1_26_port, 
        fourth_out_1_25_port, fourth_out_1_24_port, fourth_out_1_23_port, 
        fourth_out_1_22_port, fourth_out_1_21_port, fourth_out_1_20_port, 
        fourth_out_1_19_port, fourth_out_1_18_port, fourth_out_1_17_port, 
        fourth_out_1_16_port, fourth_out_1_15_port, fourth_out_1_14_port, 
        fourth_out_1_13_port, fourth_out_1_12_port, fourth_out_1_11_port, 
        fourth_out_1_10_port, fourth_out_1_9_port, fourth_out_1_8_port, 
        fourth_out_1_7_port, fourth_out_1_6_port, fourth_out_1_5_port, 
        fourth_out_1_4_port, fourth_out_1_3_port, fourth_out_1_2_port, 
        fourth_out_1_1_port, fourth_out_1_0_port}), .cout({
        fourth_cout_1_31_port, fourth_cout_1_30_port, fourth_cout_1_29_port, 
        fourth_cout_1_28_port, fourth_cout_1_27_port, fourth_cout_1_26_port, 
        fourth_cout_1_25_port, fourth_cout_1_24_port, fourth_cout_1_23_port, 
        fourth_cout_1_22_port, fourth_cout_1_21_port, fourth_cout_1_20_port, 
        fourth_cout_1_19_port, fourth_cout_1_18_port, fourth_cout_1_17_port, 
        fourth_cout_1_16_port, fourth_cout_1_15_port, fourth_cout_1_14_port, 
        fourth_cout_1_13_port, fourth_cout_1_12_port, fourth_cout_1_11_port, 
        fourth_cout_1_10_port, fourth_cout_1_9_port, fourth_cout_1_8_port, 
        fourth_cout_1_7_port, fourth_cout_1_6_port, fourth_cout_1_5_port, 
        fourth_cout_1_4_port, fourth_cout_1_3_port, fourth_cout_1_2_port, 
        fourth_cout_1_1_port, SYNOPSYS_UNCONNECTED__11}) );
  CSA_N32_2 CSA12 ( .A({fourth_out_0_31_port, fourth_out_0_30_port, 
        fourth_out_0_29_port, fourth_out_0_28_port, fourth_out_0_27_port, 
        fourth_out_0_26_port, fourth_out_0_25_port, fourth_out_0_24_port, 
        fourth_out_0_23_port, fourth_out_0_22_port, fourth_out_0_21_port, 
        fourth_out_0_20_port, fourth_out_0_19_port, fourth_out_0_18_port, 
        fourth_out_0_17_port, fourth_out_0_16_port, fourth_out_0_15_port, 
        fourth_out_0_14_port, fourth_out_0_13_port, fourth_out_0_12_port, 
        fourth_out_0_11_port, fourth_out_0_10_port, fourth_out_0_9_port, 
        fourth_out_0_8_port, fourth_out_0_7_port, fourth_out_0_6_port, 
        fourth_out_0_5_port, fourth_out_0_4_port, fourth_out_0_3_port, 
        fourth_out_0_2_port, fourth_out_0_1_port, fourth_out_0_0_port}), .B({
        fourth_cout_0_31_port, fourth_cout_0_30_port, fourth_cout_0_29_port, 
        fourth_cout_0_28_port, fourth_cout_0_27_port, fourth_cout_0_26_port, 
        fourth_cout_0_25_port, fourth_cout_0_24_port, fourth_cout_0_23_port, 
        fourth_cout_0_22_port, fourth_cout_0_21_port, fourth_cout_0_20_port, 
        fourth_cout_0_19_port, fourth_cout_0_18_port, fourth_cout_0_17_port, 
        fourth_cout_0_16_port, fourth_cout_0_15_port, fourth_cout_0_14_port, 
        fourth_cout_0_13_port, fourth_cout_0_12_port, fourth_cout_0_11_port, 
        fourth_cout_0_10_port, fourth_cout_0_9_port, fourth_cout_0_8_port, 
        fourth_cout_0_7_port, fourth_cout_0_6_port, fourth_cout_0_5_port, 
        fourth_cout_0_4_port, fourth_cout_0_3_port, fourth_cout_0_2_port, 
        fourth_cout_0_1_port, 1'b0}), .C({fourth_out_1_31_port, 
        fourth_out_1_30_port, fourth_out_1_29_port, fourth_out_1_28_port, 
        fourth_out_1_27_port, fourth_out_1_26_port, fourth_out_1_25_port, 
        fourth_out_1_24_port, fourth_out_1_23_port, fourth_out_1_22_port, 
        fourth_out_1_21_port, fourth_out_1_20_port, fourth_out_1_19_port, 
        fourth_out_1_18_port, fourth_out_1_17_port, fourth_out_1_16_port, 
        fourth_out_1_15_port, fourth_out_1_14_port, fourth_out_1_13_port, 
        fourth_out_1_12_port, fourth_out_1_11_port, fourth_out_1_10_port, 
        fourth_out_1_9_port, fourth_out_1_8_port, fourth_out_1_7_port, 
        fourth_out_1_6_port, fourth_out_1_5_port, fourth_out_1_4_port, 
        fourth_out_1_3_port, fourth_out_1_2_port, fourth_out_1_1_port, 
        fourth_out_1_0_port}), .sum_out({fifth_out_31_port, fifth_out_30_port, 
        fifth_out_29_port, fifth_out_28_port, fifth_out_27_port, 
        fifth_out_26_port, fifth_out_25_port, fifth_out_24_port, 
        fifth_out_23_port, fifth_out_22_port, fifth_out_21_port, 
        fifth_out_20_port, fifth_out_19_port, fifth_out_18_port, 
        fifth_out_17_port, fifth_out_16_port, fifth_out_15_port, 
        fifth_out_14_port, fifth_out_13_port, fifth_out_12_port, 
        fifth_out_11_port, fifth_out_10_port, fifth_out_9_port, 
        fifth_out_8_port, fifth_out_7_port, fifth_out_6_port, fifth_out_5_port, 
        fifth_out_4_port, fifth_out_3_port, fifth_out_2_port, fifth_out_1_port, 
        fifth_out_0_port}), .cout({fifth_cout_31_port, fifth_cout_30_port, 
        fifth_cout_29_port, fifth_cout_28_port, fifth_cout_27_port, 
        fifth_cout_26_port, fifth_cout_25_port, fifth_cout_24_port, 
        fifth_cout_23_port, fifth_cout_22_port, fifth_cout_21_port, 
        fifth_cout_20_port, fifth_cout_19_port, fifth_cout_18_port, 
        fifth_cout_17_port, fifth_cout_16_port, fifth_cout_15_port, 
        fifth_cout_14_port, fifth_cout_13_port, fifth_cout_12_port, 
        fifth_cout_11_port, fifth_cout_10_port, fifth_cout_9_port, 
        fifth_cout_8_port, fifth_cout_7_port, fifth_cout_6_port, 
        fifth_cout_5_port, fifth_cout_4_port, fifth_cout_3_port, 
        fifth_cout_2_port, fifth_cout_1_port, SYNOPSYS_UNCONNECTED__12}) );
  CSA_N32_1 CSA13 ( .A({fifth_out_31_port, fifth_out_30_port, 
        fifth_out_29_port, fifth_out_28_port, fifth_out_27_port, 
        fifth_out_26_port, fifth_out_25_port, fifth_out_24_port, 
        fifth_out_23_port, fifth_out_22_port, fifth_out_21_port, 
        fifth_out_20_port, fifth_out_19_port, fifth_out_18_port, 
        fifth_out_17_port, fifth_out_16_port, fifth_out_15_port, 
        fifth_out_14_port, fifth_out_13_port, fifth_out_12_port, 
        fifth_out_11_port, fifth_out_10_port, fifth_out_9_port, 
        fifth_out_8_port, fifth_out_7_port, fifth_out_6_port, fifth_out_5_port, 
        fifth_out_4_port, fifth_out_3_port, fifth_out_2_port, fifth_out_1_port, 
        fifth_out_0_port}), .B({fifth_cout_31_port, fifth_cout_30_port, 
        fifth_cout_29_port, fifth_cout_28_port, fifth_cout_27_port, 
        fifth_cout_26_port, fifth_cout_25_port, fifth_cout_24_port, 
        fifth_cout_23_port, fifth_cout_22_port, fifth_cout_21_port, 
        fifth_cout_20_port, fifth_cout_19_port, fifth_cout_18_port, 
        fifth_cout_17_port, fifth_cout_16_port, fifth_cout_15_port, 
        fifth_cout_14_port, fifth_cout_13_port, fifth_cout_12_port, 
        fifth_cout_11_port, fifth_cout_10_port, fifth_cout_9_port, 
        fifth_cout_8_port, fifth_cout_7_port, fifth_cout_6_port, 
        fifth_cout_5_port, fifth_cout_4_port, fifth_cout_3_port, 
        fifth_cout_2_port, fifth_cout_1_port, 1'b0}), .C({
        fourth_cout_1_31_port, fourth_cout_1_30_port, fourth_cout_1_29_port, 
        fourth_cout_1_28_port, fourth_cout_1_27_port, fourth_cout_1_26_port, 
        fourth_cout_1_25_port, fourth_cout_1_24_port, fourth_cout_1_23_port, 
        fourth_cout_1_22_port, fourth_cout_1_21_port, fourth_cout_1_20_port, 
        fourth_cout_1_19_port, fourth_cout_1_18_port, fourth_cout_1_17_port, 
        fourth_cout_1_16_port, fourth_cout_1_15_port, fourth_cout_1_14_port, 
        fourth_cout_1_13_port, fourth_cout_1_12_port, fourth_cout_1_11_port, 
        fourth_cout_1_10_port, fourth_cout_1_9_port, fourth_cout_1_8_port, 
        fourth_cout_1_7_port, fourth_cout_1_6_port, fourth_cout_1_5_port, 
        fourth_cout_1_4_port, fourth_cout_1_3_port, fourth_cout_1_2_port, 
        fourth_cout_1_1_port, 1'b0}), .sum_out({sixth_out_31_port, 
        sixth_out_30_port, sixth_out_29_port, sixth_out_28_port, 
        sixth_out_27_port, sixth_out_26_port, sixth_out_25_port, 
        sixth_out_24_port, sixth_out_23_port, sixth_out_22_port, 
        sixth_out_21_port, sixth_out_20_port, sixth_out_19_port, 
        sixth_out_18_port, sixth_out_17_port, sixth_out_16_port, 
        sixth_out_15_port, sixth_out_14_port, sixth_out_13_port, 
        sixth_out_12_port, sixth_out_11_port, sixth_out_10_port, 
        sixth_out_9_port, sixth_out_8_port, sixth_out_7_port, sixth_out_6_port, 
        sixth_out_5_port, sixth_out_4_port, sixth_out_3_port, sixth_out_2_port, 
        sixth_out_1_port, sixth_out_0_port}), .cout({sixth_cout_31_port, 
        sixth_cout_30_port, sixth_cout_29_port, sixth_cout_28_port, 
        sixth_cout_27_port, sixth_cout_26_port, sixth_cout_25_port, 
        sixth_cout_24_port, sixth_cout_23_port, sixth_cout_22_port, 
        sixth_cout_21_port, sixth_cout_20_port, sixth_cout_19_port, 
        sixth_cout_18_port, sixth_cout_17_port, sixth_cout_16_port, 
        sixth_cout_15_port, sixth_cout_14_port, sixth_cout_13_port, 
        sixth_cout_12_port, sixth_cout_11_port, sixth_cout_10_port, 
        sixth_cout_9_port, sixth_cout_8_port, sixth_cout_7_port, 
        sixth_cout_6_port, sixth_cout_5_port, sixth_cout_4_port, 
        sixth_cout_3_port, sixth_cout_2_port, sixth_cout_1_port, 
        SYNOPSYS_UNCONNECTED__13}) );
  P4adderN_Nbit32 P4A14 ( .A({sixth_out_31_port, sixth_out_30_port, 
        sixth_out_29_port, sixth_out_28_port, sixth_out_27_port, 
        sixth_out_26_port, sixth_out_25_port, sixth_out_24_port, 
        sixth_out_23_port, sixth_out_22_port, sixth_out_21_port, 
        sixth_out_20_port, sixth_out_19_port, sixth_out_18_port, 
        sixth_out_17_port, sixth_out_16_port, sixth_out_15_port, 
        sixth_out_14_port, sixth_out_13_port, sixth_out_12_port, 
        sixth_out_11_port, sixth_out_10_port, sixth_out_9_port, 
        sixth_out_8_port, sixth_out_7_port, sixth_out_6_port, sixth_out_5_port, 
        sixth_out_4_port, sixth_out_3_port, sixth_out_2_port, sixth_out_1_port, 
        sixth_out_0_port}), .B({sixth_cout_31_port, sixth_cout_30_port, 
        sixth_cout_29_port, sixth_cout_28_port, sixth_cout_27_port, 
        sixth_cout_26_port, sixth_cout_25_port, sixth_cout_24_port, 
        sixth_cout_23_port, sixth_cout_22_port, sixth_cout_21_port, 
        sixth_cout_20_port, sixth_cout_19_port, sixth_cout_18_port, 
        sixth_cout_17_port, sixth_cout_16_port, sixth_cout_15_port, 
        sixth_cout_14_port, sixth_cout_13_port, sixth_cout_12_port, 
        sixth_cout_11_port, sixth_cout_10_port, sixth_cout_9_port, 
        sixth_cout_8_port, sixth_cout_7_port, sixth_cout_6_port, 
        sixth_cout_5_port, sixth_cout_4_port, sixth_cout_3_port, 
        sixth_cout_2_port, sixth_cout_1_port, 1'b0}), .Cin(1'b0), .S(p) );
  BoothMulWallace_Nbit32_DW01_inc_0 add_72 ( .A({N132, N35, N36, N37, N38, N39, 
        N40, N41, N42, N43, N44, N45, N46, N47, N48, N49}), .SUM({N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50})
         );
  NOR2_X2 U4 ( .A1(n65), .A2(n68), .ZN(n420) );
  NOR2_X2 U5 ( .A1(n65), .A2(n69), .ZN(n418) );
  NOR2_X2 U6 ( .A1(n70), .A2(n65), .ZN(n411) );
  NOR2_X2 U34 ( .A1(n65), .A2(n102), .ZN(init_8_31_port) );
  AOI21_X2 U48 ( .B1(a[8]), .B2(n103), .A(n104), .ZN(n102) );
  AOI21_X2 U104 ( .B1(a[5]), .B2(n103), .A(n122), .ZN(n121) );
  AOI21_X2 U140 ( .B1(a[3]), .B2(n103), .A(n132), .ZN(n78) );
  AOI22_X2 U271 ( .A1(a[11]), .A2(n103), .B1(n158), .B2(n167), .ZN(n70) );
  AOI21_X2 U308 ( .B1(a[9]), .B2(n255), .A(n176), .ZN(n85) );
  AOI21_X2 U313 ( .B1(a[8]), .B2(n255), .A(n178), .ZN(n86) );
  AOI21_X2 U317 ( .B1(a[7]), .B2(n255), .A(n180), .ZN(n71) );
  AOI21_X2 U322 ( .B1(a[6]), .B2(n255), .A(n182), .ZN(n73) );
  AOI21_X2 U327 ( .B1(a[5]), .B2(n255), .A(n184), .ZN(n87) );
  AOI21_X2 U331 ( .B1(a[4]), .B2(n255), .A(n186), .ZN(n88) );
  AOI21_X2 U336 ( .B1(a[3]), .B2(n255), .A(n188), .ZN(n89) );
  AOI21_X2 U340 ( .B1(a[2]), .B2(n255), .A(n190), .ZN(n90) );
  AOI21_X2 U345 ( .B1(a[1]), .B2(n255), .A(n192), .ZN(n91) );
  AOI21_X2 U349 ( .B1(a[14]), .B2(n255), .A(n194), .ZN(n80) );
  AOI21_X2 U354 ( .B1(a[13]), .B2(n255), .A(n196), .ZN(n81) );
  AOI21_X2 U359 ( .B1(a[12]), .B2(n255), .A(n198), .ZN(n82) );
  AOI21_X2 U364 ( .B1(a[11]), .B2(n256), .A(n200), .ZN(n83) );
  AOI21_X2 U369 ( .B1(a[10]), .B2(n256), .A(n202), .ZN(n84) );
  AOI21_X2 U374 ( .B1(a[0]), .B2(n256), .A(n204), .ZN(n79) );
  AOI22_X2 U378 ( .A1(n100), .A2(b[0]), .B1(a[0]), .B2(n103), .ZN(n75) );
  NAND3_X1 U402 ( .A1(n97), .A2(n94), .A3(n98), .ZN(n96) );
  NAND3_X1 U403 ( .A1(n107), .A2(n252), .A3(b[8]), .ZN(n106) );
  NAND3_X1 U404 ( .A1(n100), .A2(n109), .A3(n110), .ZN(n107) );
  NAND3_X1 U405 ( .A1(n114), .A2(n109), .A3(n98), .ZN(n113) );
  NAND3_X1 U406 ( .A1(n119), .A2(n117), .A3(n98), .ZN(n118) );
  NAND3_X1 U407 ( .A1(n125), .A2(n252), .A3(b[5]), .ZN(n124) );
  NAND3_X1 U408 ( .A1(n100), .A2(n126), .A3(n127), .ZN(n125) );
  NAND3_X1 U409 ( .A1(n131), .A2(n126), .A3(n98), .ZN(n130) );
  NAND3_X1 U410 ( .A1(n135), .A2(n252), .A3(b[3]), .ZN(n134) );
  NAND3_X1 U411 ( .A1(n100), .A2(n136), .A3(n137), .ZN(n135) );
  NAND3_X1 U412 ( .A1(n141), .A2(n136), .A3(n98), .ZN(n140) );
  NAND3_X1 U413 ( .A1(n98), .A2(n147), .A3(n148), .ZN(n72) );
  NAND3_X1 U414 ( .A1(n158), .A2(n160), .A3(n98), .ZN(n165) );
  INV_X1 U2 ( .A(n154), .ZN(n153) );
  NOR2_X1 U3 ( .A1(n65), .A2(n161), .ZN(init_12_31_port) );
  OR2_X1 U7 ( .A1(n98), .A2(n103), .ZN(n252) );
  NOR2_X4 U8 ( .A1(n65), .A2(n67), .ZN(n425) );
  INV_X2 U9 ( .A(n253), .ZN(init_5_31_port) );
  NOR2_X4 U10 ( .A1(n65), .A2(n66), .ZN(n431) );
  INV_X1 U11 ( .A(n150), .ZN(n149) );
  INV_X1 U12 ( .A(n92), .ZN(n69) );
  INV_X1 U13 ( .A(n252), .ZN(n255) );
  INV_X1 U14 ( .A(n252), .ZN(n256) );
  INV_X1 U15 ( .A(n146), .ZN(n100) );
  INV_X1 U16 ( .A(n254), .ZN(n103) );
  BUF_X2 U17 ( .A(n250), .Z(n257) );
  BUF_X2 U18 ( .A(n247), .Z(n263) );
  BUF_X2 U19 ( .A(n248), .Z(n261) );
  BUF_X2 U20 ( .A(n249), .Z(n259) );
  NOR2_X1 U21 ( .A1(n98), .A2(n256), .ZN(n146) );
  BUF_X1 U22 ( .A(n250), .Z(n258) );
  BUF_X1 U23 ( .A(n249), .Z(n260) );
  BUF_X1 U24 ( .A(n248), .Z(n262) );
  INV_X1 U25 ( .A(n166), .ZN(n158) );
  NAND2_X1 U26 ( .A1(n100), .A2(n160), .ZN(n159) );
  NAND2_X1 U27 ( .A1(n100), .A2(n173), .ZN(n172) );
  BUF_X1 U28 ( .A(n247), .Z(n264) );
  INV_X1 U29 ( .A(n137), .ZN(n141) );
  INV_X1 U30 ( .A(n144), .ZN(n98) );
  NOR2_X1 U31 ( .A1(n65), .A2(n153), .ZN(init_13_31_port) );
  NOR2_X1 U32 ( .A1(n65), .A2(n72), .ZN(init_15_31_port) );
  NOR2_X1 U33 ( .A1(n65), .A2(n149), .ZN(init_14_31_port) );
  OR2_X1 U35 ( .A1(n65), .A2(n121), .ZN(n253) );
  NAND2_X1 U36 ( .A1(b[15]), .A2(N132), .ZN(n95) );
  NAND2_X1 U37 ( .A1(b[15]), .A2(N132), .ZN(n254) );
  NOR3_X1 U38 ( .A1(b[10]), .A2(b[11]), .A3(n171), .ZN(n166) );
  NOR2_X1 U39 ( .A1(n81), .A2(n72), .ZN(init_15_28_port) );
  NOR2_X1 U40 ( .A1(n82), .A2(n72), .ZN(init_15_27_port) );
  NOR2_X1 U41 ( .A1(n83), .A2(n72), .ZN(init_15_26_port) );
  NOR2_X1 U42 ( .A1(n85), .A2(n72), .ZN(init_15_24_port) );
  NOR2_X1 U43 ( .A1(n86), .A2(n72), .ZN(init_15_23_port) );
  NOR2_X1 U44 ( .A1(n71), .A2(n72), .ZN(n410) );
  NOR2_X1 U45 ( .A1(n87), .A2(n72), .ZN(init_15_20_port) );
  NOR2_X1 U46 ( .A1(n88), .A2(n72), .ZN(init_15_19_port) );
  NOR2_X1 U47 ( .A1(n89), .A2(n72), .ZN(init_15_18_port) );
  NOR2_X1 U49 ( .A1(n91), .A2(n72), .ZN(init_15_16_port) );
  NOR2_X1 U50 ( .A1(n79), .A2(n72), .ZN(init_15_15_port) );
  NOR2_X1 U51 ( .A1(n80), .A2(n72), .ZN(init_15_29_port) );
  NOR2_X1 U52 ( .A1(n84), .A2(n72), .ZN(init_15_25_port) );
  NOR2_X1 U53 ( .A1(n73), .A2(n72), .ZN(n409) );
  NOR2_X1 U54 ( .A1(n90), .A2(n72), .ZN(init_15_17_port) );
  INV_X1 U55 ( .A(n138), .ZN(n77) );
  OAI221_X1 U56 ( .B1(n139), .B2(n136), .C1(N47), .C2(n95), .A(n140), .ZN(n138) );
  AOI21_X1 U57 ( .B1(n137), .B2(n100), .A(n256), .ZN(n139) );
  INV_X1 U58 ( .A(n115), .ZN(n66) );
  OAI221_X1 U59 ( .B1(n116), .B2(n117), .C1(N43), .C2(n95), .A(n118), .ZN(n115) );
  AOI21_X1 U60 ( .B1(n120), .B2(n100), .A(n256), .ZN(n116) );
  INV_X1 U61 ( .A(n163), .ZN(n161) );
  OAI221_X1 U62 ( .B1(n164), .B2(n160), .C1(N37), .C2(n95), .A(n165), .ZN(n163) );
  AOI21_X1 U63 ( .B1(n166), .B2(n100), .A(n256), .ZN(n164) );
  INV_X1 U64 ( .A(n111), .ZN(n67) );
  OAI221_X1 U65 ( .B1(n112), .B2(n109), .C1(N42), .C2(n254), .A(n113), .ZN(
        n111) );
  AOI21_X1 U66 ( .B1(n110), .B2(n100), .A(n256), .ZN(n112) );
  INV_X1 U67 ( .A(n128), .ZN(n74) );
  OAI221_X1 U68 ( .B1(n129), .B2(n126), .C1(N45), .C2(n254), .A(n130), .ZN(
        n128) );
  AOI21_X1 U69 ( .B1(n127), .B2(n100), .A(n256), .ZN(n129) );
  NOR2_X1 U70 ( .A1(n80), .A2(n70), .ZN(init_11_25_port) );
  NOR2_X1 U71 ( .A1(n81), .A2(n70), .ZN(init_11_24_port) );
  NOR2_X1 U72 ( .A1(n82), .A2(n70), .ZN(init_11_23_port) );
  NOR2_X1 U73 ( .A1(n83), .A2(n70), .ZN(init_11_22_port) );
  NOR2_X1 U74 ( .A1(n84), .A2(n70), .ZN(init_11_21_port) );
  NOR2_X1 U75 ( .A1(n85), .A2(n70), .ZN(init_11_20_port) );
  NOR2_X1 U76 ( .A1(n86), .A2(n70), .ZN(init_11_19_port) );
  NOR2_X1 U77 ( .A1(n71), .A2(n70), .ZN(init_11_18_port) );
  NOR2_X1 U78 ( .A1(n73), .A2(n70), .ZN(init_11_17_port) );
  NOR2_X1 U79 ( .A1(n87), .A2(n70), .ZN(init_11_16_port) );
  NOR2_X1 U80 ( .A1(n88), .A2(n70), .ZN(init_11_15_port) );
  NOR2_X1 U81 ( .A1(n89), .A2(n70), .ZN(init_11_14_port) );
  NOR2_X1 U82 ( .A1(n90), .A2(n70), .ZN(init_11_13_port) );
  NOR2_X1 U83 ( .A1(n91), .A2(n70), .ZN(init_11_12_port) );
  NOR2_X1 U84 ( .A1(n79), .A2(n70), .ZN(init_11_11_port) );
  NOR2_X1 U85 ( .A1(n75), .A2(n80), .ZN(init_0_14_port) );
  NOR2_X1 U86 ( .A1(n75), .A2(n82), .ZN(init_0_12_port) );
  NOR2_X1 U87 ( .A1(n75), .A2(n83), .ZN(init_0_11_port) );
  NOR2_X1 U88 ( .A1(n75), .A2(n86), .ZN(init_0_8_port) );
  NOR2_X1 U89 ( .A1(n75), .A2(n71), .ZN(init_0_7_port) );
  NOR2_X1 U90 ( .A1(n75), .A2(n73), .ZN(init_0_6_port) );
  NOR2_X1 U91 ( .A1(n75), .A2(n88), .ZN(init_0_4_port) );
  NOR2_X1 U92 ( .A1(n75), .A2(n89), .ZN(init_0_3_port) );
  NOR2_X1 U93 ( .A1(n75), .A2(n90), .ZN(init_0_2_port) );
  NOR2_X1 U94 ( .A1(n75), .A2(n84), .ZN(init_0_10_port) );
  NOR2_X1 U95 ( .A1(n75), .A2(n81), .ZN(init_0_13_port) );
  NOR2_X1 U96 ( .A1(n75), .A2(n85), .ZN(init_0_9_port) );
  NOR2_X1 U97 ( .A1(n75), .A2(n87), .ZN(init_0_5_port) );
  NOR2_X1 U98 ( .A1(n75), .A2(n79), .ZN(init_0_0_port) );
  NOR2_X1 U99 ( .A1(n75), .A2(n91), .ZN(init_0_1_port) );
  NOR2_X1 U100 ( .A1(n80), .A2(n78), .ZN(init_3_17_port) );
  NOR2_X1 U101 ( .A1(n81), .A2(n78), .ZN(init_3_16_port) );
  NOR2_X1 U102 ( .A1(n82), .A2(n78), .ZN(init_3_15_port) );
  NOR2_X1 U103 ( .A1(n84), .A2(n78), .ZN(init_3_13_port) );
  NOR2_X1 U105 ( .A1(n85), .A2(n78), .ZN(init_3_12_port) );
  NOR2_X1 U106 ( .A1(n73), .A2(n78), .ZN(init_3_9_port) );
  NOR2_X1 U107 ( .A1(n87), .A2(n78), .ZN(init_3_8_port) );
  NOR2_X1 U108 ( .A1(n88), .A2(n78), .ZN(init_3_7_port) );
  NOR2_X1 U109 ( .A1(n90), .A2(n78), .ZN(init_3_5_port) );
  NOR2_X1 U110 ( .A1(n91), .A2(n78), .ZN(init_3_4_port) );
  NOR2_X1 U111 ( .A1(n79), .A2(n78), .ZN(init_3_3_port) );
  NOR2_X1 U112 ( .A1(n86), .A2(n78), .ZN(init_3_11_port) );
  NOR2_X1 U113 ( .A1(n83), .A2(n78), .ZN(init_3_14_port) );
  NOR2_X1 U114 ( .A1(n71), .A2(n78), .ZN(init_3_10_port) );
  NOR2_X1 U115 ( .A1(n89), .A2(n78), .ZN(init_3_6_port) );
  NOR2_X1 U116 ( .A1(n80), .A2(n121), .ZN(init_5_19_port) );
  NOR2_X1 U117 ( .A1(n82), .A2(n121), .ZN(init_5_17_port) );
  NOR2_X1 U118 ( .A1(n83), .A2(n121), .ZN(init_5_16_port) );
  NOR2_X1 U119 ( .A1(n84), .A2(n121), .ZN(init_5_15_port) );
  NOR2_X1 U120 ( .A1(n86), .A2(n121), .ZN(init_5_13_port) );
  NOR2_X1 U121 ( .A1(n71), .A2(n121), .ZN(init_5_12_port) );
  NOR2_X1 U122 ( .A1(n88), .A2(n121), .ZN(init_5_9_port) );
  NOR2_X1 U123 ( .A1(n89), .A2(n121), .ZN(init_5_8_port) );
  NOR2_X1 U124 ( .A1(n90), .A2(n121), .ZN(init_5_7_port) );
  NOR2_X1 U125 ( .A1(n79), .A2(n121), .ZN(init_5_5_port) );
  NOR2_X1 U126 ( .A1(n73), .A2(n121), .ZN(init_5_11_port) );
  NOR2_X1 U127 ( .A1(n80), .A2(n102), .ZN(init_8_22_port) );
  NOR2_X1 U128 ( .A1(n81), .A2(n102), .ZN(init_8_21_port) );
  NOR2_X1 U129 ( .A1(n82), .A2(n102), .ZN(init_8_20_port) );
  NOR2_X1 U130 ( .A1(n83), .A2(n102), .ZN(init_8_19_port) );
  NOR2_X1 U131 ( .A1(n84), .A2(n102), .ZN(init_8_18_port) );
  NOR2_X1 U132 ( .A1(n81), .A2(n121), .ZN(init_5_18_port) );
  NOR2_X1 U133 ( .A1(n85), .A2(n102), .ZN(init_8_17_port) );
  NOR2_X1 U134 ( .A1(n86), .A2(n102), .ZN(init_8_16_port) );
  NOR2_X1 U135 ( .A1(n71), .A2(n102), .ZN(init_8_15_port) );
  NOR2_X1 U136 ( .A1(n73), .A2(n102), .ZN(init_8_14_port) );
  NOR2_X1 U137 ( .A1(n85), .A2(n121), .ZN(init_5_14_port) );
  NOR2_X1 U138 ( .A1(n87), .A2(n102), .ZN(init_8_13_port) );
  NOR2_X1 U139 ( .A1(n90), .A2(n102), .ZN(init_8_10_port) );
  NOR2_X1 U141 ( .A1(n87), .A2(n121), .ZN(init_5_10_port) );
  NOR2_X1 U142 ( .A1(n91), .A2(n102), .ZN(init_8_9_port) );
  NOR2_X1 U143 ( .A1(n79), .A2(n102), .ZN(init_8_8_port) );
  NOR2_X1 U144 ( .A1(n91), .A2(n121), .ZN(init_5_6_port) );
  NOR2_X1 U145 ( .A1(n88), .A2(n102), .ZN(init_8_12_port) );
  NOR2_X1 U146 ( .A1(n89), .A2(n102), .ZN(init_8_11_port) );
  NOR2_X1 U147 ( .A1(n80), .A2(n69), .ZN(init_9_23_port) );
  NOR2_X1 U148 ( .A1(n81), .A2(n69), .ZN(init_9_22_port) );
  NOR2_X1 U149 ( .A1(n82), .A2(n69), .ZN(init_9_21_port) );
  NOR2_X1 U150 ( .A1(n83), .A2(n69), .ZN(init_9_20_port) );
  NOR2_X1 U151 ( .A1(n84), .A2(n69), .ZN(init_9_19_port) );
  NOR2_X1 U152 ( .A1(n80), .A2(n66), .ZN(init_6_20_port) );
  NOR2_X1 U153 ( .A1(n81), .A2(n66), .ZN(init_6_19_port) );
  NOR2_X1 U154 ( .A1(n85), .A2(n69), .ZN(init_9_18_port) );
  NOR2_X1 U155 ( .A1(n82), .A2(n66), .ZN(init_6_18_port) );
  NOR2_X1 U156 ( .A1(n86), .A2(n69), .ZN(init_9_17_port) );
  NOR2_X1 U157 ( .A1(n83), .A2(n66), .ZN(init_6_17_port) );
  NOR2_X1 U158 ( .A1(n71), .A2(n69), .ZN(init_9_16_port) );
  NOR2_X1 U159 ( .A1(n73), .A2(n69), .ZN(init_9_15_port) );
  NOR2_X1 U160 ( .A1(n84), .A2(n66), .ZN(init_6_16_port) );
  NOR2_X1 U161 ( .A1(n85), .A2(n66), .ZN(init_6_15_port) );
  NOR2_X1 U162 ( .A1(n87), .A2(n69), .ZN(init_9_14_port) );
  NOR2_X1 U163 ( .A1(n86), .A2(n66), .ZN(init_6_14_port) );
  NOR2_X1 U164 ( .A1(n88), .A2(n69), .ZN(init_9_13_port) );
  NOR2_X1 U165 ( .A1(n71), .A2(n66), .ZN(init_6_13_port) );
  NOR2_X1 U166 ( .A1(n91), .A2(n69), .ZN(init_9_10_port) );
  NOR2_X1 U167 ( .A1(n88), .A2(n66), .ZN(init_6_10_port) );
  NOR2_X1 U168 ( .A1(n79), .A2(n69), .ZN(init_9_9_port) );
  NOR2_X1 U169 ( .A1(n89), .A2(n66), .ZN(init_6_9_port) );
  NOR2_X1 U170 ( .A1(n90), .A2(n66), .ZN(init_6_8_port) );
  NOR2_X1 U171 ( .A1(n91), .A2(n66), .ZN(init_6_7_port) );
  NOR2_X1 U172 ( .A1(n79), .A2(n66), .ZN(init_6_6_port) );
  NOR2_X1 U173 ( .A1(n89), .A2(n69), .ZN(init_9_12_port) );
  NOR2_X1 U174 ( .A1(n73), .A2(n66), .ZN(init_6_12_port) );
  NOR2_X1 U175 ( .A1(n90), .A2(n69), .ZN(init_9_11_port) );
  NOR2_X1 U176 ( .A1(n87), .A2(n66), .ZN(init_6_11_port) );
  NOR2_X1 U177 ( .A1(n80), .A2(n161), .ZN(init_12_26_port) );
  NOR2_X1 U178 ( .A1(n81), .A2(n161), .ZN(init_12_25_port) );
  NOR2_X1 U179 ( .A1(n82), .A2(n161), .ZN(init_12_24_port) );
  NOR2_X1 U180 ( .A1(n83), .A2(n161), .ZN(init_12_23_port) );
  NOR2_X1 U181 ( .A1(n84), .A2(n161), .ZN(init_12_22_port) );
  NOR2_X1 U182 ( .A1(n85), .A2(n161), .ZN(init_12_21_port) );
  NOR2_X1 U183 ( .A1(n86), .A2(n161), .ZN(init_12_20_port) );
  NOR2_X1 U184 ( .A1(n71), .A2(n161), .ZN(init_12_19_port) );
  NOR2_X1 U185 ( .A1(n73), .A2(n161), .ZN(init_12_18_port) );
  NOR2_X1 U186 ( .A1(n87), .A2(n161), .ZN(init_12_17_port) );
  NOR2_X1 U187 ( .A1(n88), .A2(n161), .ZN(init_12_16_port) );
  NOR2_X1 U188 ( .A1(n89), .A2(n161), .ZN(init_12_15_port) );
  NOR2_X1 U189 ( .A1(n90), .A2(n161), .ZN(init_12_14_port) );
  NOR2_X1 U190 ( .A1(n91), .A2(n161), .ZN(init_12_13_port) );
  NOR2_X1 U191 ( .A1(n79), .A2(n161), .ZN(init_12_12_port) );
  NOR2_X1 U192 ( .A1(n80), .A2(n77), .ZN(init_2_16_port) );
  NOR2_X1 U193 ( .A1(n81), .A2(n77), .ZN(init_2_15_port) );
  NOR2_X1 U194 ( .A1(n82), .A2(n77), .ZN(init_2_14_port) );
  NOR2_X1 U195 ( .A1(n84), .A2(n77), .ZN(init_2_12_port) );
  NOR2_X1 U196 ( .A1(n85), .A2(n77), .ZN(init_2_11_port) );
  NOR2_X1 U197 ( .A1(n73), .A2(n77), .ZN(init_2_8_port) );
  NOR2_X1 U198 ( .A1(n87), .A2(n77), .ZN(init_2_7_port) );
  NOR2_X1 U199 ( .A1(n88), .A2(n77), .ZN(init_2_6_port) );
  NOR2_X1 U200 ( .A1(n90), .A2(n77), .ZN(init_2_4_port) );
  NOR2_X1 U201 ( .A1(n91), .A2(n77), .ZN(init_2_3_port) );
  NOR2_X1 U202 ( .A1(n79), .A2(n77), .ZN(init_2_2_port) );
  NOR2_X1 U203 ( .A1(n86), .A2(n77), .ZN(init_2_10_port) );
  NOR2_X1 U204 ( .A1(n83), .A2(n77), .ZN(init_2_13_port) );
  NOR2_X1 U205 ( .A1(n71), .A2(n77), .ZN(init_2_9_port) );
  NOR2_X1 U206 ( .A1(n89), .A2(n77), .ZN(init_2_5_port) );
  NOR2_X1 U207 ( .A1(n81), .A2(n149), .ZN(init_14_27_port) );
  NOR2_X1 U208 ( .A1(n82), .A2(n149), .ZN(init_14_26_port) );
  NOR2_X1 U209 ( .A1(n83), .A2(n149), .ZN(init_14_25_port) );
  NOR2_X1 U210 ( .A1(n84), .A2(n149), .ZN(init_14_24_port) );
  NOR2_X1 U211 ( .A1(n85), .A2(n149), .ZN(init_14_23_port) );
  NOR2_X1 U212 ( .A1(n86), .A2(n149), .ZN(init_14_22_port) );
  NOR2_X1 U213 ( .A1(n71), .A2(n149), .ZN(init_14_21_port) );
  NOR2_X1 U214 ( .A1(n73), .A2(n149), .ZN(init_14_20_port) );
  NOR2_X1 U215 ( .A1(n87), .A2(n149), .ZN(init_14_19_port) );
  NOR2_X1 U216 ( .A1(n88), .A2(n149), .ZN(init_14_18_port) );
  NOR2_X1 U217 ( .A1(n89), .A2(n149), .ZN(init_14_17_port) );
  NOR2_X1 U218 ( .A1(n90), .A2(n149), .ZN(init_14_16_port) );
  NOR2_X1 U219 ( .A1(n91), .A2(n149), .ZN(init_14_15_port) );
  NOR2_X1 U220 ( .A1(n79), .A2(n149), .ZN(init_14_14_port) );
  NOR2_X1 U221 ( .A1(n80), .A2(n149), .ZN(init_14_28_port) );
  NOR2_X1 U222 ( .A1(n80), .A2(n76), .ZN(init_1_15_port) );
  NOR2_X1 U223 ( .A1(n81), .A2(n76), .ZN(init_1_14_port) );
  NOR2_X1 U224 ( .A1(n83), .A2(n76), .ZN(init_1_12_port) );
  NOR2_X1 U225 ( .A1(n84), .A2(n76), .ZN(init_1_11_port) );
  NOR2_X1 U226 ( .A1(n71), .A2(n76), .ZN(init_1_8_port) );
  NOR2_X1 U227 ( .A1(n73), .A2(n76), .ZN(init_1_7_port) );
  NOR2_X1 U228 ( .A1(n87), .A2(n76), .ZN(init_1_6_port) );
  NOR2_X1 U229 ( .A1(n89), .A2(n76), .ZN(init_1_4_port) );
  NOR2_X1 U230 ( .A1(n90), .A2(n76), .ZN(init_1_3_port) );
  NOR2_X1 U231 ( .A1(n91), .A2(n76), .ZN(init_1_2_port) );
  NOR2_X1 U232 ( .A1(n85), .A2(n76), .ZN(init_1_10_port) );
  NOR2_X1 U233 ( .A1(n82), .A2(n76), .ZN(init_1_13_port) );
  NOR2_X1 U234 ( .A1(n86), .A2(n76), .ZN(init_1_9_port) );
  NOR2_X1 U235 ( .A1(n88), .A2(n76), .ZN(init_1_5_port) );
  NOR2_X1 U236 ( .A1(n81), .A2(n74), .ZN(init_4_17_port) );
  NOR2_X1 U237 ( .A1(n82), .A2(n74), .ZN(init_4_16_port) );
  NOR2_X1 U238 ( .A1(n83), .A2(n74), .ZN(init_4_15_port) );
  NOR2_X1 U239 ( .A1(n85), .A2(n74), .ZN(init_4_13_port) );
  NOR2_X1 U240 ( .A1(n86), .A2(n74), .ZN(init_4_12_port) );
  NOR2_X1 U241 ( .A1(n87), .A2(n74), .ZN(init_4_9_port) );
  NOR2_X1 U242 ( .A1(n88), .A2(n74), .ZN(init_4_8_port) );
  NOR2_X1 U243 ( .A1(n89), .A2(n74), .ZN(init_4_7_port) );
  NOR2_X1 U244 ( .A1(n91), .A2(n74), .ZN(init_4_5_port) );
  NOR2_X1 U245 ( .A1(n79), .A2(n74), .ZN(init_4_4_port) );
  NOR2_X1 U246 ( .A1(n79), .A2(n76), .ZN(init_1_1_port) );
  NOR2_X1 U247 ( .A1(n71), .A2(n74), .ZN(init_4_11_port) );
  NOR2_X1 U248 ( .A1(n80), .A2(n68), .ZN(init_10_24_port) );
  NOR2_X1 U249 ( .A1(n81), .A2(n68), .ZN(init_10_23_port) );
  NOR2_X1 U250 ( .A1(n82), .A2(n68), .ZN(init_10_22_port) );
  NOR2_X1 U251 ( .A1(n83), .A2(n68), .ZN(init_10_21_port) );
  NOR2_X1 U252 ( .A1(n80), .A2(n67), .ZN(init_7_21_port) );
  NOR2_X1 U253 ( .A1(n84), .A2(n68), .ZN(init_10_20_port) );
  NOR2_X1 U254 ( .A1(n85), .A2(n68), .ZN(init_10_19_port) );
  NOR2_X1 U255 ( .A1(n81), .A2(n67), .ZN(init_7_20_port) );
  NOR2_X1 U256 ( .A1(n82), .A2(n67), .ZN(init_7_19_port) );
  NOR2_X1 U257 ( .A1(n86), .A2(n68), .ZN(init_10_18_port) );
  NOR2_X1 U258 ( .A1(n83), .A2(n67), .ZN(init_7_18_port) );
  NOR2_X1 U259 ( .A1(n80), .A2(n74), .ZN(init_4_18_port) );
  NOR2_X1 U260 ( .A1(n71), .A2(n68), .ZN(init_10_17_port) );
  NOR2_X1 U261 ( .A1(n84), .A2(n67), .ZN(init_7_17_port) );
  NOR2_X1 U262 ( .A1(n73), .A2(n68), .ZN(init_10_16_port) );
  NOR2_X1 U263 ( .A1(n87), .A2(n68), .ZN(init_10_15_port) );
  NOR2_X1 U264 ( .A1(n85), .A2(n67), .ZN(init_7_16_port) );
  NOR2_X1 U265 ( .A1(n86), .A2(n67), .ZN(init_7_15_port) );
  NOR2_X1 U266 ( .A1(n88), .A2(n68), .ZN(init_10_14_port) );
  NOR2_X1 U267 ( .A1(n71), .A2(n67), .ZN(init_7_14_port) );
  NOR2_X1 U268 ( .A1(n84), .A2(n74), .ZN(init_4_14_port) );
  NOR2_X1 U269 ( .A1(n89), .A2(n68), .ZN(init_10_13_port) );
  NOR2_X1 U270 ( .A1(n73), .A2(n67), .ZN(init_7_13_port) );
  NOR2_X1 U272 ( .A1(n79), .A2(n68), .ZN(init_10_10_port) );
  NOR2_X1 U273 ( .A1(n89), .A2(n67), .ZN(init_7_10_port) );
  NOR2_X1 U274 ( .A1(n73), .A2(n74), .ZN(init_4_10_port) );
  NOR2_X1 U275 ( .A1(n90), .A2(n67), .ZN(init_7_9_port) );
  NOR2_X1 U276 ( .A1(n91), .A2(n67), .ZN(init_7_8_port) );
  NOR2_X1 U277 ( .A1(n79), .A2(n67), .ZN(init_7_7_port) );
  NOR2_X1 U278 ( .A1(n90), .A2(n74), .ZN(init_4_6_port) );
  NOR2_X1 U279 ( .A1(n90), .A2(n68), .ZN(init_10_12_port) );
  NOR2_X1 U280 ( .A1(n87), .A2(n67), .ZN(init_7_12_port) );
  NOR2_X1 U281 ( .A1(n91), .A2(n68), .ZN(init_10_11_port) );
  NOR2_X1 U282 ( .A1(n88), .A2(n67), .ZN(init_7_11_port) );
  NOR2_X1 U283 ( .A1(n80), .A2(n153), .ZN(init_13_27_port) );
  NOR2_X1 U284 ( .A1(n81), .A2(n153), .ZN(init_13_26_port) );
  NOR2_X1 U285 ( .A1(n82), .A2(n153), .ZN(init_13_25_port) );
  NOR2_X1 U286 ( .A1(n83), .A2(n153), .ZN(init_13_24_port) );
  NOR2_X1 U287 ( .A1(n84), .A2(n153), .ZN(init_13_23_port) );
  NOR2_X1 U288 ( .A1(n85), .A2(n153), .ZN(init_13_22_port) );
  NOR2_X1 U289 ( .A1(n86), .A2(n153), .ZN(init_13_21_port) );
  NOR2_X1 U290 ( .A1(n71), .A2(n153), .ZN(init_13_20_port) );
  NOR2_X1 U291 ( .A1(n73), .A2(n153), .ZN(init_13_19_port) );
  NOR2_X1 U292 ( .A1(n87), .A2(n153), .ZN(init_13_18_port) );
  NOR2_X1 U293 ( .A1(n88), .A2(n153), .ZN(init_13_17_port) );
  NOR2_X1 U294 ( .A1(n89), .A2(n153), .ZN(init_13_16_port) );
  NOR2_X1 U295 ( .A1(n90), .A2(n153), .ZN(init_13_15_port) );
  NOR2_X1 U296 ( .A1(n91), .A2(n153), .ZN(init_13_14_port) );
  NOR2_X1 U297 ( .A1(n79), .A2(n153), .ZN(init_13_13_port) );
  NOR2_X1 U298 ( .A1(n75), .A2(n65), .ZN(n250) );
  NOR2_X1 U299 ( .A1(n65), .A2(n78), .ZN(n247) );
  NOR2_X1 U300 ( .A1(b[1]), .A2(b[0]), .ZN(n137) );
  NOR2_X1 U301 ( .A1(n65), .A2(n77), .ZN(n248) );
  NOR2_X1 U302 ( .A1(n65), .A2(n76), .ZN(n249) );
  INV_X1 U303 ( .A(b[0]), .ZN(n145) );
  INV_X1 U304 ( .A(b[12]), .ZN(n160) );
  NOR2_X1 U305 ( .A1(n74), .A2(n65), .ZN(n443) );
  INV_X1 U306 ( .A(n127), .ZN(n131) );
  INV_X1 U307 ( .A(b[10]), .ZN(n173) );
  INV_X1 U309 ( .A(n99), .ZN(n97) );
  INV_X1 U310 ( .A(n120), .ZN(n119) );
  INV_X1 U311 ( .A(b[11]), .ZN(n168) );
  INV_X1 U312 ( .A(n110), .ZN(n114) );
  OAI22_X1 U314 ( .A1(n168), .A2(n169), .B1(n144), .B2(b[11]), .ZN(n167) );
  INV_X1 U315 ( .A(n170), .ZN(n169) );
  OAI21_X1 U316 ( .B1(n171), .B2(n172), .A(n252), .ZN(n170) );
  INV_X1 U318 ( .A(n133), .ZN(n132) );
  OAI211_X1 U319 ( .C1(b[3]), .C2(n98), .A(n134), .B(n131), .ZN(n133) );
  INV_X1 U320 ( .A(n105), .ZN(n104) );
  OAI211_X1 U321 ( .C1(b[8]), .C2(n98), .A(n106), .B(n97), .ZN(n105) );
  INV_X1 U323 ( .A(n123), .ZN(n122) );
  OAI211_X1 U324 ( .C1(b[5]), .C2(n98), .A(n124), .B(n119), .ZN(n123) );
  OAI22_X1 U325 ( .A1(n195), .A2(n144), .B1(n147), .B2(n254), .ZN(n194) );
  INV_X1 U326 ( .A(N64), .ZN(n195) );
  OAI22_X1 U328 ( .A1(n199), .A2(n144), .B1(n160), .B2(n254), .ZN(n198) );
  INV_X1 U329 ( .A(N62), .ZN(n199) );
  INV_X1 U330 ( .A(n179), .ZN(n178) );
  AOI22_X1 U332 ( .A1(N58), .A2(n98), .B1(b[8]), .B2(n103), .ZN(n179) );
  OAI22_X1 U333 ( .A1(n181), .A2(n144), .B1(n109), .B2(n95), .ZN(n180) );
  INV_X1 U334 ( .A(N57), .ZN(n181) );
  OAI22_X1 U335 ( .A1(n183), .A2(n144), .B1(n117), .B2(n254), .ZN(n182) );
  INV_X1 U337 ( .A(N56), .ZN(n183) );
  OAI22_X1 U338 ( .A1(n187), .A2(n144), .B1(n254), .B2(n126), .ZN(n186) );
  INV_X1 U339 ( .A(N54), .ZN(n187) );
  INV_X1 U341 ( .A(n189), .ZN(n188) );
  AOI22_X1 U342 ( .A1(N53), .A2(n98), .B1(b[3]), .B2(n103), .ZN(n189) );
  OAI22_X1 U343 ( .A1(n191), .A2(n144), .B1(n136), .B2(n95), .ZN(n190) );
  INV_X1 U344 ( .A(N52), .ZN(n191) );
  OAI22_X1 U346 ( .A1(n197), .A2(n144), .B1(n157), .B2(n95), .ZN(n196) );
  INV_X1 U347 ( .A(N63), .ZN(n197) );
  OAI22_X1 U348 ( .A1(n177), .A2(n144), .B1(n94), .B2(n254), .ZN(n176) );
  INV_X1 U350 ( .A(N59), .ZN(n177) );
  INV_X1 U351 ( .A(n185), .ZN(n184) );
  AOI22_X1 U352 ( .A1(N55), .A2(n98), .B1(b[5]), .B2(n103), .ZN(n185) );
  INV_X1 U353 ( .A(n193), .ZN(n192) );
  AOI22_X1 U355 ( .A1(N51), .A2(n98), .B1(b[1]), .B2(n103), .ZN(n193) );
  OAI22_X1 U356 ( .A1(n201), .A2(n144), .B1(n168), .B2(n95), .ZN(n200) );
  INV_X1 U357 ( .A(N61), .ZN(n201) );
  OAI22_X1 U358 ( .A1(n203), .A2(n144), .B1(n173), .B2(n254), .ZN(n202) );
  INV_X1 U360 ( .A(N60), .ZN(n203) );
  OAI22_X1 U361 ( .A1(n205), .A2(n144), .B1(n145), .B2(n95), .ZN(n204) );
  INV_X1 U362 ( .A(N50), .ZN(n205) );
  OAI22_X1 U363 ( .A1(N36), .A2(n95), .B1(n148), .B2(n155), .ZN(n154) );
  AOI22_X1 U365 ( .A1(b[13]), .A2(n156), .B1(n98), .B2(n157), .ZN(n155) );
  OAI21_X1 U366 ( .B1(n158), .B2(n159), .A(n252), .ZN(n156) );
  NAND2_X1 U367 ( .A1(b[15]), .A2(a[15]), .ZN(n144) );
  NOR3_X1 U368 ( .A1(b[12]), .A2(b[13]), .A3(n158), .ZN(n148) );
  NOR3_X1 U370 ( .A1(b[7]), .A2(b[8]), .A3(n114), .ZN(n99) );
  NOR3_X1 U371 ( .A1(b[2]), .A2(b[3]), .A3(n141), .ZN(n127) );
  NOR3_X1 U372 ( .A1(b[4]), .A2(b[5]), .A3(n131), .ZN(n120) );
  OAI21_X1 U373 ( .B1(n146), .B2(b[0]), .A(n252), .ZN(n142) );
  NOR3_X1 U375 ( .A1(n144), .A2(b[1]), .A3(n145), .ZN(n143) );
  AND3_X1 U376 ( .A1(n171), .A2(n173), .A3(n98), .ZN(n175) );
  OAI21_X1 U377 ( .B1(n171), .B2(n146), .A(n252), .ZN(n174) );
  AND2_X1 U379 ( .A1(N65), .A2(n98), .ZN(n162) );
  OAI221_X1 U380 ( .B1(n93), .B2(n94), .C1(N40), .C2(n95), .A(n96), .ZN(n92)
         );
  AOI21_X1 U381 ( .B1(n99), .B2(n100), .A(n256), .ZN(n93) );
  OAI221_X1 U382 ( .B1(n151), .B2(n147), .C1(N35), .C2(n254), .A(n152), .ZN(
        n150) );
  OR3_X1 U383 ( .A1(n148), .A2(b[14]), .A3(n144), .ZN(n152) );
  AOI21_X1 U384 ( .B1(n148), .B2(n100), .A(n256), .ZN(n151) );
  NOR2_X1 U385 ( .A1(n119), .A2(b[6]), .ZN(n110) );
  NAND2_X1 U386 ( .A1(n99), .A2(n94), .ZN(n171) );
  INV_X1 U387 ( .A(a[6]), .ZN(N43) );
  INV_X1 U388 ( .A(a[14]), .ZN(N35) );
  INV_X1 U389 ( .A(a[12]), .ZN(N37) );
  INV_X1 U390 ( .A(a[2]), .ZN(N47) );
  INV_X1 U391 ( .A(b[13]), .ZN(n157) );
  INV_X1 U392 ( .A(b[4]), .ZN(n126) );
  INV_X1 U393 ( .A(b[2]), .ZN(n136) );
  INV_X1 U394 ( .A(b[7]), .ZN(n109) );
  INV_X1 U395 ( .A(a[15]), .ZN(N132) );
  INV_X1 U396 ( .A(a[9]), .ZN(N40) );
  INV_X1 U397 ( .A(a[7]), .ZN(N42) );
  INV_X1 U398 ( .A(a[13]), .ZN(N36) );
  INV_X1 U399 ( .A(b[14]), .ZN(n147) );
  INV_X1 U400 ( .A(a[4]), .ZN(N45) );
  INV_X1 U401 ( .A(b[6]), .ZN(n117) );
  INV_X1 U415 ( .A(a[3]), .ZN(N46) );
  INV_X1 U416 ( .A(a[8]), .ZN(N41) );
  INV_X1 U417 ( .A(a[5]), .ZN(N44) );
  INV_X1 U418 ( .A(a[10]), .ZN(N39) );
  INV_X1 U419 ( .A(a[1]), .ZN(N48) );
  INV_X1 U420 ( .A(a[0]), .ZN(N49) );
  INV_X1 U421 ( .A(a[11]), .ZN(N38) );
  INV_X1 U422 ( .A(b[9]), .ZN(n94) );
  AOI221_X4 U423 ( .B1(n174), .B2(b[10]), .C1(a[10]), .C2(n103), .A(n175), 
        .ZN(n68) );
  AOI211_X4 U424 ( .C1(a[15]), .C2(n256), .A(n103), .B(n162), .ZN(n65) );
  AOI221_X4 U425 ( .B1(n142), .B2(b[1]), .C1(a[1]), .C2(n103), .A(n143), .ZN(
        n76) );
  CLKBUF_X1 U426 ( .A(n443), .Z(n265) );
  CLKBUF_X1 U427 ( .A(n443), .Z(n266) );
endmodule


module mux21N_N32_4 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;

  tri   S;

  MUX21_288 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_287 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_286 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_285 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_284 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
  MUX21_283 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(S), .Y(U[5]) );
  MUX21_282 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(S), .Y(U[6]) );
  MUX21_281 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(S), .Y(U[7]) );
  MUX21_280 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(S), .Y(U[8]) );
  MUX21_279 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(S), .Y(U[9]) );
  MUX21_278 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(S), .Y(U[10]) );
  MUX21_277 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(S), .Y(U[11]) );
  MUX21_276 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(S), .Y(U[12]) );
  MUX21_275 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(S), .Y(U[13]) );
  MUX21_274 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(S), .Y(U[14]) );
  MUX21_273 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(S), .Y(U[15]) );
  MUX21_272 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(S), .Y(U[16]) );
  MUX21_271 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(S), .Y(U[17]) );
  MUX21_270 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(S), .Y(U[18]) );
  MUX21_269 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(S), .Y(U[19]) );
  MUX21_268 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(S), .Y(U[20]) );
  MUX21_267 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(S), .Y(U[21]) );
  MUX21_266 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(S), .Y(U[22]) );
  MUX21_265 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(S), .Y(U[23]) );
  MUX21_264 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(S), .Y(U[24]) );
  MUX21_263 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(S), .Y(U[25]) );
  MUX21_262 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(S), .Y(U[26]) );
  MUX21_261 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(S), .Y(U[27]) );
  MUX21_260 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(S), .Y(U[28]) );
  MUX21_259 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(S), .Y(U[29]) );
  MUX21_258 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(S), .Y(U[30]) );
  MUX21_257 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(S), .Y(U[31]) );
endmodule


module mux21N_N32_5 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   net399734, n37, n38, n39, n40, n41, n42;
  assign net399734 = S;

  MUX21_320 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n42), .Y(U[0]) );
  MUX21_319 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n38), .Y(U[1]) );
  MUX21_318 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n42), .Y(U[2]) );
  MUX21_317 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n39), .Y(U[3]) );
  MUX21_316 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n38), .Y(U[4]) );
  MUX21_315 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n37), .Y(U[5]) );
  MUX21_314 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n38), .Y(U[6]) );
  MUX21_313 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n42), .Y(U[7]) );
  MUX21_312 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n38), .Y(U[8]) );
  MUX21_311 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n42), .Y(U[9]) );
  MUX21_310 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n38), .Y(U[10]) );
  MUX21_309 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n42), .Y(U[11]) );
  MUX21_308 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n38), .Y(U[12]) );
  MUX21_307 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n42), .Y(U[13]) );
  MUX21_306 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n40), .Y(U[14]) );
  MUX21_305 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n42), .Y(U[15]) );
  MUX21_304 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n40), .Y(U[16]) );
  MUX21_303 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n40), .Y(U[17]) );
  MUX21_302 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n38), .Y(U[18]) );
  MUX21_301 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n40), .Y(U[19]) );
  MUX21_300 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n37), .Y(U[20]) );
  MUX21_299 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n39), .Y(U[21]) );
  MUX21_298 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n40), .Y(U[22]) );
  MUX21_297 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n39), .Y(U[23]) );
  MUX21_296 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n40), .Y(U[24]) );
  MUX21_295 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n40), .Y(U[25]) );
  MUX21_294 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n37), .Y(U[26]) );
  MUX21_293 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n40), .Y(U[27]) );
  MUX21_292 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n40), .Y(U[28]) );
  MUX21_291 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n40), .Y(U[29]) );
  MUX21_290 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n40), .Y(U[30]) );
  MUX21_289 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n40), .Y(U[31]) );
  BUF_X2 U1 ( .A(n41), .Z(n39) );
  CLKBUF_X3 U2 ( .A(net399734), .Z(n42) );
  BUF_X1 U3 ( .A(net399734), .Z(n41) );
  BUF_X4 U4 ( .A(net399734), .Z(n40) );
  BUF_X1 U5 ( .A(n41), .Z(n37) );
  CLKBUF_X3 U6 ( .A(n41), .Z(n38) );
endmodule


module mux21N_N32_6 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   net397599, n20, n21, n22, n23;
  assign net397599 = S;

  MUX21_352 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n23), .Y(U[0]) );
  MUX21_351 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n21), .Y(U[1]) );
  MUX21_350 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n22), .Y(U[2]) );
  MUX21_349 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n23), .Y(U[3]) );
  MUX21_348 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n21), .Y(U[4]) );
  MUX21_347 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n21), .Y(U[5]) );
  MUX21_346 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n21), .Y(U[6]) );
  MUX21_345 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n22), .Y(U[7]) );
  MUX21_344 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n21), .Y(U[8]) );
  MUX21_343 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n22), .Y(U[9]) );
  MUX21_342 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n22), .Y(U[10]) );
  MUX21_341 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n22), .Y(U[11]) );
  MUX21_340 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n21), .Y(U[12]) );
  MUX21_339 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n22), .Y(U[13]) );
  MUX21_338 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n21), .Y(U[14]) );
  MUX21_337 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n23), .Y(U[15]) );
  MUX21_336 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n21), .Y(U[16]) );
  MUX21_335 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n23), .Y(U[17]) );
  MUX21_334 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n22), .Y(U[18]) );
  MUX21_333 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n23), .Y(U[19]) );
  MUX21_332 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n22), .Y(U[20]) );
  MUX21_331 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n23), .Y(U[21]) );
  MUX21_330 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n21), .Y(U[22]) );
  MUX21_329 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n22), .Y(U[23]) );
  MUX21_328 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n21), .Y(U[24]) );
  MUX21_327 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n20), .Y(U[25]) );
  MUX21_326 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n22), .Y(U[26]) );
  MUX21_325 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n22), .Y(U[27]) );
  MUX21_324 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n20), .Y(U[28]) );
  MUX21_323 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n20), .Y(U[29]) );
  MUX21_322 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n21), .Y(U[30]) );
  MUX21_321 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n20), .Y(U[31]) );
  CLKBUF_X3 U1 ( .A(net397599), .Z(n22) );
  CLKBUF_X2 U2 ( .A(net397599), .Z(n21) );
  BUF_X2 U3 ( .A(n23), .Z(n20) );
  CLKBUF_X2 U4 ( .A(net397599), .Z(n23) );
endmodule


module MUX21_479 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_486 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_491 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_493 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_494 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_497 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_498 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_499 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_501 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_502 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module CarrySumN_Nbit32_2 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  CSBlockN_Nbit4_16 CSN_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  CSBlockN_Nbit4_15 CSN_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  CSBlockN_Nbit4_14 CSN_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8])
         );
  CSBlockN_Nbit4_13 CSN_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  CSBlockN_Nbit4_12 CSN_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  CSBlockN_Nbit4_11 CSN_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  CSBlockN_Nbit4_10 CSN_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  CSBlockN_Nbit4_9 CSN_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(S[31:28]) );
endmodule


module SparseTreeCarryGenN_Nbit32_2 ( A, B, Cin, Cout );
  input [31:0] A;
  input [31:0] B;
  output [8:0] Cout;
  input Cin;
  wire   Cin, propcin, gencin, \gen[4][28] , \gen[4][32] , \gen[3][16] ,
         \gen[3][24] , \gen[3][32] , \gen[2][8] , \gen[2][12] , \gen[2][16] ,
         \gen[2][20] , \gen[2][24] , \gen[2][28] , \gen[2][32] , \gen[1][2] ,
         \gen[1][4] , \gen[1][6] , \gen[1][8] , \gen[1][10] , \gen[1][12] ,
         \gen[1][14] , \gen[1][16] , \gen[1][18] , \gen[1][20] , \gen[1][22] ,
         \gen[1][24] , \gen[1][26] , \gen[1][28] , \gen[1][30] , \gen[1][32] ,
         \gen[0][1] , \gen[0][2] , \gen[0][3] , \gen[0][4] , \gen[0][5] ,
         \gen[0][6] , \gen[0][7] , \gen[0][8] , \gen[0][9] , \gen[0][10] ,
         \gen[0][11] , \gen[0][12] , \gen[0][13] , \gen[0][14] , \gen[0][15] ,
         \gen[0][16] , \gen[0][17] , \gen[0][18] , \gen[0][19] , \gen[0][20] ,
         \gen[0][21] , \gen[0][22] , \gen[0][23] , \gen[0][24] , \gen[0][25] ,
         \gen[0][26] , \gen[0][27] , \gen[0][28] , \gen[0][29] , \gen[0][30] ,
         \gen[0][31] , \gen[0][32] , \prop[4][28] , \prop[4][32] ,
         \prop[3][16] , \prop[3][24] , \prop[3][32] , \prop[2][8] ,
         \prop[2][12] , \prop[2][16] , \prop[2][20] , \prop[2][24] ,
         \prop[2][28] , \prop[2][32] , \prop[1][4] , \prop[1][6] ,
         \prop[1][8] , \prop[1][10] , \prop[1][12] , \prop[1][14] ,
         \prop[1][16] , \prop[1][18] , \prop[1][20] , \prop[1][22] ,
         \prop[1][24] , \prop[1][26] , \prop[1][28] , \prop[1][30] ,
         \prop[1][32] , \prop[0][2] , \prop[0][3] , \prop[0][4] , \prop[0][5] ,
         \prop[0][6] , \prop[0][7] , \prop[0][8] , \prop[0][9] , \prop[0][10] ,
         \prop[0][11] , \prop[0][12] , \prop[0][13] , \prop[0][14] ,
         \prop[0][15] , \prop[0][16] , \prop[0][17] , \prop[0][18] ,
         \prop[0][19] , \prop[0][20] , \prop[0][21] , \prop[0][22] ,
         \prop[0][23] , \prop[0][24] , \prop[0][25] , \prop[0][26] ,
         \prop[0][27] , \prop[0][28] , \prop[0][29] , \prop[0][30] ,
         \prop[0][31] , \prop[0][32] , n2;
  assign Cout[0] = Cin;

  PGblock_96 Cinprop_0_1 ( .A(A[0]), .B(B[0]), .G(gencin), .P(propcin) );
  PGblock_95 PGB_0_2 ( .A(A[1]), .B(B[1]), .G(\gen[0][2] ), .P(\prop[0][2] )
         );
  PGblock_94 PGB_0_3 ( .A(A[2]), .B(B[2]), .G(\gen[0][3] ), .P(\prop[0][3] )
         );
  PGblock_93 PGB_0_4 ( .A(A[3]), .B(B[3]), .G(\gen[0][4] ), .P(\prop[0][4] )
         );
  PGblock_92 PGB_0_5 ( .A(A[4]), .B(B[4]), .G(\gen[0][5] ), .P(\prop[0][5] )
         );
  PGblock_91 PGB_0_6 ( .A(A[5]), .B(B[5]), .G(\gen[0][6] ), .P(\prop[0][6] )
         );
  PGblock_90 PGB_0_7 ( .A(A[6]), .B(B[6]), .G(\gen[0][7] ), .P(\prop[0][7] )
         );
  PGblock_89 PGB_0_8 ( .A(A[7]), .B(B[7]), .G(\gen[0][8] ), .P(\prop[0][8] )
         );
  PGblock_88 PGB_0_9 ( .A(A[8]), .B(B[8]), .G(\gen[0][9] ), .P(\prop[0][9] )
         );
  PGblock_87 PGB_0_10 ( .A(A[9]), .B(B[9]), .G(\gen[0][10] ), .P(\prop[0][10] ) );
  PGblock_86 PGB_0_11 ( .A(A[10]), .B(B[10]), .G(\gen[0][11] ), .P(
        \prop[0][11] ) );
  PGblock_85 PGB_0_12 ( .A(A[11]), .B(B[11]), .G(\gen[0][12] ), .P(
        \prop[0][12] ) );
  PGblock_84 PGB_0_13 ( .A(A[12]), .B(B[12]), .G(\gen[0][13] ), .P(
        \prop[0][13] ) );
  PGblock_83 PGB_0_14 ( .A(A[13]), .B(B[13]), .G(\gen[0][14] ), .P(
        \prop[0][14] ) );
  PGblock_82 PGB_0_15 ( .A(A[14]), .B(B[14]), .G(\gen[0][15] ), .P(
        \prop[0][15] ) );
  PGblock_81 PGB_0_16 ( .A(A[15]), .B(B[15]), .G(\gen[0][16] ), .P(
        \prop[0][16] ) );
  PGblock_80 PGB_0_17 ( .A(A[16]), .B(B[16]), .G(\gen[0][17] ), .P(
        \prop[0][17] ) );
  PGblock_79 PGB_0_18 ( .A(A[17]), .B(B[17]), .G(\gen[0][18] ), .P(
        \prop[0][18] ) );
  PGblock_78 PGB_0_19 ( .A(A[18]), .B(B[18]), .G(\gen[0][19] ), .P(
        \prop[0][19] ) );
  PGblock_77 PGB_0_20 ( .A(A[19]), .B(B[19]), .G(\gen[0][20] ), .P(
        \prop[0][20] ) );
  PGblock_76 PGB_0_21 ( .A(A[20]), .B(B[20]), .G(\gen[0][21] ), .P(
        \prop[0][21] ) );
  PGblock_75 PGB_0_22 ( .A(A[21]), .B(B[21]), .G(\gen[0][22] ), .P(
        \prop[0][22] ) );
  PGblock_74 PGB_0_23 ( .A(A[22]), .B(B[22]), .G(\gen[0][23] ), .P(
        \prop[0][23] ) );
  PGblock_73 PGB_0_24 ( .A(A[23]), .B(B[23]), .G(\gen[0][24] ), .P(
        \prop[0][24] ) );
  PGblock_72 PGB_0_25 ( .A(A[24]), .B(B[24]), .G(\gen[0][25] ), .P(
        \prop[0][25] ) );
  PGblock_71 PGB_0_26 ( .A(A[25]), .B(B[25]), .G(\gen[0][26] ), .P(
        \prop[0][26] ) );
  PGblock_70 PGB_0_27 ( .A(A[26]), .B(B[26]), .G(\gen[0][27] ), .P(
        \prop[0][27] ) );
  PGblock_69 PGB_0_28 ( .A(A[27]), .B(B[27]), .G(\gen[0][28] ), .P(
        \prop[0][28] ) );
  PGblock_68 PGB_0_29 ( .A(A[28]), .B(B[28]), .G(\gen[0][29] ), .P(
        \prop[0][29] ) );
  PGblock_67 PGB_0_30 ( .A(A[29]), .B(B[29]), .G(\gen[0][30] ), .P(
        \prop[0][30] ) );
  PGblock_66 PGB_0_31 ( .A(A[30]), .B(B[30]), .G(\gen[0][31] ), .P(
        \prop[0][31] ) );
  PGblock_65 PGB_0_32 ( .A(A[31]), .B(B[31]), .G(\gen[0][32] ), .P(
        \prop[0][32] ) );
  G_27 G1_2_1_1 ( .G1(\gen[0][2] ), .P1(\prop[0][2] ), .G2(\gen[0][1] ), 
        .Gout(\gen[1][2] ) );
  PG_81 PG1_2_1_2 ( .G1(\gen[0][4] ), .P1(\prop[0][4] ), .G2(\gen[0][3] ), 
        .P2(\prop[0][3] ), .Gout(\gen[1][4] ), .Pout(\prop[1][4] ) );
  PG_80 PG1_2_1_3 ( .G1(\gen[0][6] ), .P1(\prop[0][6] ), .G2(\gen[0][5] ), 
        .P2(\prop[0][5] ), .Gout(\gen[1][6] ), .Pout(\prop[1][6] ) );
  PG_79 PG1_2_1_4 ( .G1(\gen[0][8] ), .P1(\prop[0][8] ), .G2(\gen[0][7] ), 
        .P2(\prop[0][7] ), .Gout(\gen[1][8] ), .Pout(\prop[1][8] ) );
  PG_78 PG1_2_1_5 ( .G1(\gen[0][10] ), .P1(\prop[0][10] ), .G2(\gen[0][9] ), 
        .P2(\prop[0][9] ), .Gout(\gen[1][10] ), .Pout(\prop[1][10] ) );
  PG_77 PG1_2_1_6 ( .G1(\gen[0][12] ), .P1(\prop[0][12] ), .G2(\gen[0][11] ), 
        .P2(\prop[0][11] ), .Gout(\gen[1][12] ), .Pout(\prop[1][12] ) );
  PG_76 PG1_2_1_7 ( .G1(\gen[0][14] ), .P1(\prop[0][14] ), .G2(\gen[0][13] ), 
        .P2(\prop[0][13] ), .Gout(\gen[1][14] ), .Pout(\prop[1][14] ) );
  PG_75 PG1_2_1_8 ( .G1(\gen[0][16] ), .P1(\prop[0][16] ), .G2(\gen[0][15] ), 
        .P2(\prop[0][15] ), .Gout(\gen[1][16] ), .Pout(\prop[1][16] ) );
  PG_74 PG1_2_1_9 ( .G1(\gen[0][18] ), .P1(\prop[0][18] ), .G2(\gen[0][17] ), 
        .P2(\prop[0][17] ), .Gout(\gen[1][18] ), .Pout(\prop[1][18] ) );
  PG_73 PG1_2_1_10 ( .G1(\gen[0][20] ), .P1(\prop[0][20] ), .G2(\gen[0][19] ), 
        .P2(\prop[0][19] ), .Gout(\gen[1][20] ), .Pout(\prop[1][20] ) );
  PG_72 PG1_2_1_11 ( .G1(\gen[0][22] ), .P1(\prop[0][22] ), .G2(\gen[0][21] ), 
        .P2(\prop[0][21] ), .Gout(\gen[1][22] ), .Pout(\prop[1][22] ) );
  PG_71 PG1_2_1_12 ( .G1(\gen[0][24] ), .P1(\prop[0][24] ), .G2(\gen[0][23] ), 
        .P2(\prop[0][23] ), .Gout(\gen[1][24] ), .Pout(\prop[1][24] ) );
  PG_70 PG1_2_1_13 ( .G1(\gen[0][26] ), .P1(\prop[0][26] ), .G2(\gen[0][25] ), 
        .P2(\prop[0][25] ), .Gout(\gen[1][26] ), .Pout(\prop[1][26] ) );
  PG_69 PG1_2_1_14 ( .G1(\gen[0][28] ), .P1(\prop[0][28] ), .G2(\gen[0][27] ), 
        .P2(\prop[0][27] ), .Gout(\gen[1][28] ), .Pout(\prop[1][28] ) );
  PG_68 PG1_2_1_15 ( .G1(\gen[0][30] ), .P1(\prop[0][30] ), .G2(\gen[0][29] ), 
        .P2(\prop[0][29] ), .Gout(\gen[1][30] ), .Pout(\prop[1][30] ) );
  PG_67 PG1_2_1_16 ( .G1(\gen[0][32] ), .P1(\prop[0][32] ), .G2(\gen[0][31] ), 
        .P2(\prop[0][31] ), .Gout(\gen[1][32] ), .Pout(\prop[1][32] ) );
  G_26 G1_2_2_1 ( .G1(\gen[1][4] ), .P1(\prop[1][4] ), .G2(\gen[1][2] ), 
        .Gout(Cout[1]) );
  PG_66 PG1_2_2_2 ( .G1(\gen[1][8] ), .P1(\prop[1][8] ), .G2(\gen[1][6] ), 
        .P2(\prop[1][6] ), .Gout(\gen[2][8] ), .Pout(\prop[2][8] ) );
  PG_65 PG1_2_2_3 ( .G1(\gen[1][12] ), .P1(\prop[1][12] ), .G2(\gen[1][10] ), 
        .P2(\prop[1][10] ), .Gout(\gen[2][12] ), .Pout(\prop[2][12] ) );
  PG_64 PG1_2_2_4 ( .G1(\gen[1][16] ), .P1(\prop[1][16] ), .G2(\gen[1][14] ), 
        .P2(\prop[1][14] ), .Gout(\gen[2][16] ), .Pout(\prop[2][16] ) );
  PG_63 PG1_2_2_5 ( .G1(\gen[1][20] ), .P1(\prop[1][20] ), .G2(\gen[1][18] ), 
        .P2(\prop[1][18] ), .Gout(\gen[2][20] ), .Pout(\prop[2][20] ) );
  PG_62 PG1_2_2_6 ( .G1(\gen[1][24] ), .P1(\prop[1][24] ), .G2(\gen[1][22] ), 
        .P2(\prop[1][22] ), .Gout(\gen[2][24] ), .Pout(\prop[2][24] ) );
  PG_61 PG1_2_2_7 ( .G1(\gen[1][28] ), .P1(\prop[1][28] ), .G2(\gen[1][26] ), 
        .P2(\prop[1][26] ), .Gout(\gen[2][28] ), .Pout(\prop[2][28] ) );
  PG_60 PG1_2_2_8 ( .G1(\gen[1][32] ), .P1(\prop[1][32] ), .G2(\gen[1][30] ), 
        .P2(\prop[1][30] ), .Gout(\gen[2][32] ), .Pout(\prop[2][32] ) );
  G_25 G3_3_2 ( .G1(\gen[2][8] ), .P1(\prop[2][8] ), .G2(Cout[1]), .Gout(
        Cout[2]) );
  PG_59 PG3_3_4 ( .G1(\gen[2][16] ), .P1(\prop[2][16] ), .G2(\gen[2][12] ), 
        .P2(\prop[2][12] ), .Gout(\gen[3][16] ), .Pout(\prop[3][16] ) );
  PG_58 PG3_3_6 ( .G1(\gen[2][24] ), .P1(\prop[2][24] ), .G2(\gen[2][20] ), 
        .P2(\prop[2][20] ), .Gout(\gen[3][24] ), .Pout(\prop[3][24] ) );
  PG_57 PG3_3_8 ( .G1(\gen[2][32] ), .P1(\prop[2][32] ), .G2(\gen[2][28] ), 
        .P2(\prop[2][28] ), .Gout(\gen[3][32] ), .Pout(\prop[3][32] ) );
  G_24 G3_E_4_2 ( .G1(\gen[2][12] ), .P1(\prop[2][12] ), .G2(Cout[2]), .Gout(
        Cout[3]) );
  G_23 G3_E_4_3 ( .G1(\gen[3][16] ), .P1(\prop[3][16] ), .G2(Cout[2]), .Gout(
        Cout[4]) );
  PG_56 PG3_E_4_6 ( .G1(\gen[2][28] ), .P1(\prop[2][28] ), .G2(\gen[3][24] ), 
        .P2(\prop[3][24] ), .Gout(\gen[4][28] ), .Pout(\prop[4][28] ) );
  PG_55 PG3_E_4_7 ( .G1(\gen[3][32] ), .P1(\prop[3][32] ), .G2(\gen[3][24] ), 
        .P2(\prop[3][24] ), .Gout(\gen[4][32] ), .Pout(\prop[4][32] ) );
  G_22 G3_E_5_4 ( .G1(\gen[2][20] ), .P1(\prop[2][20] ), .G2(Cout[4]), .Gout(
        Cout[5]) );
  G_21 G3_E_5_5 ( .G1(\gen[3][24] ), .P1(\prop[3][24] ), .G2(Cout[4]), .Gout(
        Cout[6]) );
  G_20 G3_E_5_6 ( .G1(\gen[4][28] ), .P1(\prop[4][28] ), .G2(Cout[4]), .Gout(
        Cout[7]) );
  G_19 G3_E_5_7 ( .G1(\gen[4][32] ), .P1(\prop[4][32] ), .G2(Cout[4]), .Gout(
        Cout[8]) );
  INV_X1 U1 ( .A(n2), .ZN(\gen[0][1] ) );
  AOI21_X1 U2 ( .B1(propcin), .B2(Cin), .A(gencin), .ZN(n2) );
endmodule


module mux21N_N5_33 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;

  tri   S;

  MUX21_357 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_356 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_355 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_354 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_353 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_34 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;

  tri   S;

  MUX21_362 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_361 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_360 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_359 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_358 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_35 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;

  tri   S;

  MUX21_367 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_366 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_365 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_364 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_363 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module MUX21_572 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_573 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_574 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_575 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_576 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module FD_EN_372 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n3) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
endmodule


module FD_EN_373 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n3) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
endmodule


module FD_EN_375 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n3) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
endmodule


module FD_EN_376 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n3) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
endmodule


module FD_EN_377 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n3) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
endmodule


module FD_EN_378 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n3) );
  NOR2_X1 U4 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U5 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
endmodule


module MUX21_648 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n10;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n10) );
endmodule


module FD_EN_428 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module FD_EN_429 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module FD_EN_430 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module FD_EN_431 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module MUX21_701 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module MUX21_702 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(S), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(Y) );
  AOI22_X1 U3 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
endmodule


module MUX21_703 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;
  tri   S;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module CarrySumN_Nbit32_0 ( A, B, Ci, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Ci;
  output [31:0] S;


  CSBlockN_Nbit4_0 CSN_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(Ci[0]), .S(S[3:0]) );
  CSBlockN_Nbit4_23 CSN_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(Ci[1]), .S(S[7:4]) );
  CSBlockN_Nbit4_22 CSN_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(Ci[2]), .S(S[11:8])
         );
  CSBlockN_Nbit4_21 CSN_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(Ci[3]), .S(
        S[15:12]) );
  CSBlockN_Nbit4_20 CSN_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(Ci[4]), .S(
        S[19:16]) );
  CSBlockN_Nbit4_19 CSN_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(Ci[5]), .S(
        S[23:20]) );
  CSBlockN_Nbit4_18 CSN_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(Ci[6]), .S(
        S[27:24]) );
  CSBlockN_Nbit4_17 CSN_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(Ci[7]), .S(
        S[31:28]) );
endmodule


module SparseTreeCarryGenN_Nbit32_0 ( A, B, Cin, Cout );
  input [31:0] A;
  input [31:0] B;
  output [8:0] Cout;
  input Cin;
  wire   Cin, propcin, gencin, \gen[4][28] , \gen[4][32] , \gen[3][16] ,
         \gen[3][24] , \gen[3][32] , \gen[2][8] , \gen[2][12] , \gen[2][16] ,
         \gen[2][20] , \gen[2][24] , \gen[2][28] , \gen[2][32] , \gen[1][2] ,
         \gen[1][4] , \gen[1][6] , \gen[1][8] , \gen[1][10] , \gen[1][12] ,
         \gen[1][14] , \gen[1][16] , \gen[1][18] , \gen[1][20] , \gen[1][22] ,
         \gen[1][24] , \gen[1][26] , \gen[1][28] , \gen[1][30] , \gen[1][32] ,
         \gen[0][1] , \gen[0][2] , \gen[0][3] , \gen[0][4] , \gen[0][5] ,
         \gen[0][6] , \gen[0][7] , \gen[0][8] , \gen[0][9] , \gen[0][10] ,
         \gen[0][11] , \gen[0][12] , \gen[0][13] , \gen[0][14] , \gen[0][15] ,
         \gen[0][16] , \gen[0][17] , \gen[0][18] , \gen[0][19] , \gen[0][20] ,
         \gen[0][21] , \gen[0][22] , \gen[0][23] , \gen[0][24] , \gen[0][25] ,
         \gen[0][26] , \gen[0][27] , \gen[0][28] , \gen[0][29] , \gen[0][30] ,
         \gen[0][31] , \gen[0][32] , \prop[4][28] , \prop[4][32] ,
         \prop[3][16] , \prop[3][24] , \prop[3][32] , \prop[2][8] ,
         \prop[2][12] , \prop[2][16] , \prop[2][20] , \prop[2][24] ,
         \prop[2][28] , \prop[2][32] , \prop[1][4] , \prop[1][6] ,
         \prop[1][8] , \prop[1][10] , \prop[1][12] , \prop[1][14] ,
         \prop[1][16] , \prop[1][18] , \prop[1][20] , \prop[1][22] ,
         \prop[1][24] , \prop[1][26] , \prop[1][28] , \prop[1][30] ,
         \prop[1][32] , \prop[0][2] , \prop[0][3] , \prop[0][4] , \prop[0][5] ,
         \prop[0][6] , \prop[0][7] , \prop[0][8] , \prop[0][9] , \prop[0][10] ,
         \prop[0][11] , \prop[0][12] , \prop[0][13] , \prop[0][14] ,
         \prop[0][15] , \prop[0][16] , \prop[0][17] , \prop[0][18] ,
         \prop[0][19] , \prop[0][20] , \prop[0][21] , \prop[0][22] ,
         \prop[0][23] , \prop[0][24] , \prop[0][25] , \prop[0][26] ,
         \prop[0][27] , \prop[0][28] , \prop[0][29] , \prop[0][30] ,
         \prop[0][31] , \prop[0][32] , n2;
  assign Cout[0] = Cin;

  PGblock_32 Cinprop_0_1 ( .A(A[0]), .B(B[0]), .G(gencin), .P(propcin) );
  PGblock_127 PGB_0_2 ( .A(A[1]), .B(B[1]), .G(\gen[0][2] ), .P(\prop[0][2] )
         );
  PGblock_126 PGB_0_3 ( .A(A[2]), .B(B[2]), .G(\gen[0][3] ), .P(\prop[0][3] )
         );
  PGblock_125 PGB_0_4 ( .A(A[3]), .B(B[3]), .G(\gen[0][4] ), .P(\prop[0][4] )
         );
  PGblock_124 PGB_0_5 ( .A(A[4]), .B(B[4]), .G(\gen[0][5] ), .P(\prop[0][5] )
         );
  PGblock_123 PGB_0_6 ( .A(A[5]), .B(B[5]), .G(\gen[0][6] ), .P(\prop[0][6] )
         );
  PGblock_122 PGB_0_7 ( .A(A[6]), .B(B[6]), .G(\gen[0][7] ), .P(\prop[0][7] )
         );
  PGblock_121 PGB_0_8 ( .A(A[7]), .B(B[7]), .G(\gen[0][8] ), .P(\prop[0][8] )
         );
  PGblock_120 PGB_0_9 ( .A(A[8]), .B(B[8]), .G(\gen[0][9] ), .P(\prop[0][9] )
         );
  PGblock_119 PGB_0_10 ( .A(A[9]), .B(B[9]), .G(\gen[0][10] ), .P(
        \prop[0][10] ) );
  PGblock_118 PGB_0_11 ( .A(A[10]), .B(B[10]), .G(\gen[0][11] ), .P(
        \prop[0][11] ) );
  PGblock_117 PGB_0_12 ( .A(A[11]), .B(B[11]), .G(\gen[0][12] ), .P(
        \prop[0][12] ) );
  PGblock_116 PGB_0_13 ( .A(A[12]), .B(B[12]), .G(\gen[0][13] ), .P(
        \prop[0][13] ) );
  PGblock_115 PGB_0_14 ( .A(A[13]), .B(B[13]), .G(\gen[0][14] ), .P(
        \prop[0][14] ) );
  PGblock_114 PGB_0_15 ( .A(A[14]), .B(B[14]), .G(\gen[0][15] ), .P(
        \prop[0][15] ) );
  PGblock_113 PGB_0_16 ( .A(A[15]), .B(B[15]), .G(\gen[0][16] ), .P(
        \prop[0][16] ) );
  PGblock_112 PGB_0_17 ( .A(A[16]), .B(B[16]), .G(\gen[0][17] ), .P(
        \prop[0][17] ) );
  PGblock_111 PGB_0_18 ( .A(A[17]), .B(B[17]), .G(\gen[0][18] ), .P(
        \prop[0][18] ) );
  PGblock_110 PGB_0_19 ( .A(A[18]), .B(B[18]), .G(\gen[0][19] ), .P(
        \prop[0][19] ) );
  PGblock_109 PGB_0_20 ( .A(A[19]), .B(B[19]), .G(\gen[0][20] ), .P(
        \prop[0][20] ) );
  PGblock_108 PGB_0_21 ( .A(A[20]), .B(B[20]), .G(\gen[0][21] ), .P(
        \prop[0][21] ) );
  PGblock_107 PGB_0_22 ( .A(A[21]), .B(B[21]), .G(\gen[0][22] ), .P(
        \prop[0][22] ) );
  PGblock_106 PGB_0_23 ( .A(A[22]), .B(B[22]), .G(\gen[0][23] ), .P(
        \prop[0][23] ) );
  PGblock_105 PGB_0_24 ( .A(A[23]), .B(B[23]), .G(\gen[0][24] ), .P(
        \prop[0][24] ) );
  PGblock_104 PGB_0_25 ( .A(A[24]), .B(B[24]), .G(\gen[0][25] ), .P(
        \prop[0][25] ) );
  PGblock_103 PGB_0_26 ( .A(A[25]), .B(B[25]), .G(\gen[0][26] ), .P(
        \prop[0][26] ) );
  PGblock_102 PGB_0_27 ( .A(A[26]), .B(B[26]), .G(\gen[0][27] ), .P(
        \prop[0][27] ) );
  PGblock_101 PGB_0_28 ( .A(A[27]), .B(B[27]), .G(\gen[0][28] ), .P(
        \prop[0][28] ) );
  PGblock_100 PGB_0_29 ( .A(A[28]), .B(B[28]), .G(\gen[0][29] ), .P(
        \prop[0][29] ) );
  PGblock_99 PGB_0_30 ( .A(A[29]), .B(B[29]), .G(\gen[0][30] ), .P(
        \prop[0][30] ) );
  PGblock_98 PGB_0_31 ( .A(A[30]), .B(B[30]), .G(\gen[0][31] ), .P(
        \prop[0][31] ) );
  PGblock_97 PGB_0_32 ( .A(A[31]), .B(B[31]), .G(\gen[0][32] ), .P(
        \prop[0][32] ) );
  G_9 G1_2_1_1 ( .G1(\gen[0][2] ), .P1(\prop[0][2] ), .G2(\gen[0][1] ), .Gout(
        \gen[1][2] ) );
  PG_27 PG1_2_1_2 ( .G1(\gen[0][4] ), .P1(\prop[0][4] ), .G2(\gen[0][3] ), 
        .P2(\prop[0][3] ), .Gout(\gen[1][4] ), .Pout(\prop[1][4] ) );
  PG_107 PG1_2_1_3 ( .G1(\gen[0][6] ), .P1(\prop[0][6] ), .G2(\gen[0][5] ), 
        .P2(\prop[0][5] ), .Gout(\gen[1][6] ), .Pout(\prop[1][6] ) );
  PG_106 PG1_2_1_4 ( .G1(\gen[0][8] ), .P1(\prop[0][8] ), .G2(\gen[0][7] ), 
        .P2(\prop[0][7] ), .Gout(\gen[1][8] ), .Pout(\prop[1][8] ) );
  PG_105 PG1_2_1_5 ( .G1(\gen[0][10] ), .P1(\prop[0][10] ), .G2(\gen[0][9] ), 
        .P2(\prop[0][9] ), .Gout(\gen[1][10] ), .Pout(\prop[1][10] ) );
  PG_104 PG1_2_1_6 ( .G1(\gen[0][12] ), .P1(\prop[0][12] ), .G2(\gen[0][11] ), 
        .P2(\prop[0][11] ), .Gout(\gen[1][12] ), .Pout(\prop[1][12] ) );
  PG_103 PG1_2_1_7 ( .G1(\gen[0][14] ), .P1(\prop[0][14] ), .G2(\gen[0][13] ), 
        .P2(\prop[0][13] ), .Gout(\gen[1][14] ), .Pout(\prop[1][14] ) );
  PG_102 PG1_2_1_8 ( .G1(\gen[0][16] ), .P1(\prop[0][16] ), .G2(\gen[0][15] ), 
        .P2(\prop[0][15] ), .Gout(\gen[1][16] ), .Pout(\prop[1][16] ) );
  PG_101 PG1_2_1_9 ( .G1(\gen[0][18] ), .P1(\prop[0][18] ), .G2(\gen[0][17] ), 
        .P2(\prop[0][17] ), .Gout(\gen[1][18] ), .Pout(\prop[1][18] ) );
  PG_100 PG1_2_1_10 ( .G1(\gen[0][20] ), .P1(\prop[0][20] ), .G2(\gen[0][19] ), 
        .P2(\prop[0][19] ), .Gout(\gen[1][20] ), .Pout(\prop[1][20] ) );
  PG_99 PG1_2_1_11 ( .G1(\gen[0][22] ), .P1(\prop[0][22] ), .G2(\gen[0][21] ), 
        .P2(\prop[0][21] ), .Gout(\gen[1][22] ), .Pout(\prop[1][22] ) );
  PG_98 PG1_2_1_12 ( .G1(\gen[0][24] ), .P1(\prop[0][24] ), .G2(\gen[0][23] ), 
        .P2(\prop[0][23] ), .Gout(\gen[1][24] ), .Pout(\prop[1][24] ) );
  PG_97 PG1_2_1_13 ( .G1(\gen[0][26] ), .P1(\prop[0][26] ), .G2(\gen[0][25] ), 
        .P2(\prop[0][25] ), .Gout(\gen[1][26] ), .Pout(\prop[1][26] ) );
  PG_96 PG1_2_1_14 ( .G1(\gen[0][28] ), .P1(\prop[0][28] ), .G2(\gen[0][27] ), 
        .P2(\prop[0][27] ), .Gout(\gen[1][28] ), .Pout(\prop[1][28] ) );
  PG_95 PG1_2_1_15 ( .G1(\gen[0][30] ), .P1(\prop[0][30] ), .G2(\gen[0][29] ), 
        .P2(\prop[0][29] ), .Gout(\gen[1][30] ), .Pout(\prop[1][30] ) );
  PG_94 PG1_2_1_16 ( .G1(\gen[0][32] ), .P1(\prop[0][32] ), .G2(\gen[0][31] ), 
        .P2(\prop[0][31] ), .Gout(\gen[1][32] ), .Pout(\prop[1][32] ) );
  G_35 G1_2_2_1 ( .G1(\gen[1][4] ), .P1(\prop[1][4] ), .G2(\gen[1][2] ), 
        .Gout(Cout[1]) );
  PG_93 PG1_2_2_2 ( .G1(\gen[1][8] ), .P1(\prop[1][8] ), .G2(\gen[1][6] ), 
        .P2(\prop[1][6] ), .Gout(\gen[2][8] ), .Pout(\prop[2][8] ) );
  PG_92 PG1_2_2_3 ( .G1(\gen[1][12] ), .P1(\prop[1][12] ), .G2(\gen[1][10] ), 
        .P2(\prop[1][10] ), .Gout(\gen[2][12] ), .Pout(\prop[2][12] ) );
  PG_91 PG1_2_2_4 ( .G1(\gen[1][16] ), .P1(\prop[1][16] ), .G2(\gen[1][14] ), 
        .P2(\prop[1][14] ), .Gout(\gen[2][16] ), .Pout(\prop[2][16] ) );
  PG_90 PG1_2_2_5 ( .G1(\gen[1][20] ), .P1(\prop[1][20] ), .G2(\gen[1][18] ), 
        .P2(\prop[1][18] ), .Gout(\gen[2][20] ), .Pout(\prop[2][20] ) );
  PG_89 PG1_2_2_6 ( .G1(\gen[1][24] ), .P1(\prop[1][24] ), .G2(\gen[1][22] ), 
        .P2(\prop[1][22] ), .Gout(\gen[2][24] ), .Pout(\prop[2][24] ) );
  PG_88 PG1_2_2_7 ( .G1(\gen[1][28] ), .P1(\prop[1][28] ), .G2(\gen[1][26] ), 
        .P2(\prop[1][26] ), .Gout(\gen[2][28] ), .Pout(\prop[2][28] ) );
  PG_87 PG1_2_2_8 ( .G1(\gen[1][32] ), .P1(\prop[1][32] ), .G2(\gen[1][30] ), 
        .P2(\prop[1][30] ), .Gout(\gen[2][32] ), .Pout(\prop[2][32] ) );
  G_34 G3_3_2 ( .G1(\gen[2][8] ), .P1(\prop[2][8] ), .G2(Cout[1]), .Gout(
        Cout[2]) );
  PG_86 PG3_3_4 ( .G1(\gen[2][16] ), .P1(\prop[2][16] ), .G2(\gen[2][12] ), 
        .P2(\prop[2][12] ), .Gout(\gen[3][16] ), .Pout(\prop[3][16] ) );
  PG_85 PG3_3_6 ( .G1(\gen[2][24] ), .P1(\prop[2][24] ), .G2(\gen[2][20] ), 
        .P2(\prop[2][20] ), .Gout(\gen[3][24] ), .Pout(\prop[3][24] ) );
  PG_84 PG3_3_8 ( .G1(\gen[2][32] ), .P1(\prop[2][32] ), .G2(\gen[2][28] ), 
        .P2(\prop[2][28] ), .Gout(\gen[3][32] ), .Pout(\prop[3][32] ) );
  G_33 G3_E_4_2 ( .G1(\gen[2][12] ), .P1(\prop[2][12] ), .G2(Cout[2]), .Gout(
        Cout[3]) );
  G_32 G3_E_4_3 ( .G1(\gen[3][16] ), .P1(\prop[3][16] ), .G2(Cout[2]), .Gout(
        Cout[4]) );
  PG_83 PG3_E_4_6 ( .G1(\gen[2][28] ), .P1(\prop[2][28] ), .G2(\gen[3][24] ), 
        .P2(\prop[3][24] ), .Gout(\gen[4][28] ), .Pout(\prop[4][28] ) );
  PG_82 PG3_E_4_7 ( .G1(\gen[3][32] ), .P1(\prop[3][32] ), .G2(\gen[3][24] ), 
        .P2(\prop[3][24] ), .Gout(\gen[4][32] ), .Pout(\prop[4][32] ) );
  G_31 G3_E_5_4 ( .G1(\gen[2][20] ), .P1(\prop[2][20] ), .G2(Cout[4]), .Gout(
        Cout[5]) );
  G_30 G3_E_5_5 ( .G1(\gen[3][24] ), .P1(\prop[3][24] ), .G2(Cout[4]), .Gout(
        Cout[6]) );
  G_29 G3_E_5_6 ( .G1(\gen[4][28] ), .P1(\prop[4][28] ), .G2(Cout[4]), .Gout(
        Cout[7]) );
  G_28 G3_E_5_7 ( .G1(\gen[4][32] ), .P1(\prop[4][32] ), .G2(Cout[4]), .Gout(
        Cout[8]) );
  INV_X1 U1 ( .A(n2), .ZN(\gen[0][1] ) );
  AOI21_X1 U2 ( .B1(propcin), .B2(Cin), .A(gencin), .ZN(n2) );
endmodule


module MUX21_735 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n15;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n15) );
endmodule


module MUX21_767 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n14;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n14), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n14) );
endmodule


module MUX21_792 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n16;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n16), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n16) );
endmodule


module MUX21_793 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n15;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n15), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n15) );
endmodule


module MUX21_794 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n14;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n14), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n14) );
endmodule


module MUX21_795 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n13;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n13), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n13) );
endmodule


module MUX21_796 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n12;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n12), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n12) );
endmodule


module MUX21_797 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n11;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n11), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n11) );
endmodule


module MUX21_798 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n10;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n10), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n10) );
endmodule


module MUX21_799 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n9;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n9), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n9) );
endmodule


module mux41N_Nbit32_1 ( in3, in2, in1, in0, sel, Y );
  input [31:0] in3;
  input [31:0] in2;
  input [31:0] in1;
  input [31:0] in0;
  input [1:0] sel;
  output [31:0] Y;
  wire   \outmux[2][31] , \outmux[2][30] , \outmux[2][29] , \outmux[2][28] ,
         \outmux[2][27] , \outmux[2][26] , \outmux[2][25] , \outmux[2][24] ,
         \outmux[2][23] , \outmux[2][22] , \outmux[2][21] , \outmux[2][20] ,
         \outmux[2][19] , \outmux[2][18] , \outmux[2][17] , \outmux[2][16] ,
         \outmux[2][15] , \outmux[2][14] , \outmux[2][13] , \outmux[2][12] ,
         \outmux[2][11] , \outmux[2][10] , \outmux[2][9] , \outmux[2][8] ,
         \outmux[2][7] , \outmux[2][6] , \outmux[2][5] , \outmux[2][4] ,
         \outmux[2][3] , \outmux[2][2] , \outmux[2][1] , \outmux[2][0] ,
         \outmux[1][31] , \outmux[1][30] , \outmux[1][29] , \outmux[1][28] ,
         \outmux[1][27] , \outmux[1][26] , \outmux[1][25] , \outmux[1][24] ,
         \outmux[1][23] , \outmux[1][22] , \outmux[1][21] , \outmux[1][20] ,
         \outmux[1][19] , \outmux[1][18] , \outmux[1][17] , \outmux[1][16] ,
         \outmux[1][15] , \outmux[1][14] , \outmux[1][13] , \outmux[1][12] ,
         \outmux[1][11] , \outmux[1][10] , \outmux[1][9] , \outmux[1][8] ,
         \outmux[1][7] , \outmux[1][6] , \outmux[1][5] , \outmux[1][4] ,
         \outmux[1][3] , \outmux[1][2] , \outmux[1][1] , \outmux[1][0] ;

  mux21N_N32_3 row1_1 ( .in1(in1), .in0(in0), .S(sel[0]), .U({\outmux[1][31] , 
        \outmux[1][30] , \outmux[1][29] , \outmux[1][28] , \outmux[1][27] , 
        \outmux[1][26] , \outmux[1][25] , \outmux[1][24] , \outmux[1][23] , 
        \outmux[1][22] , \outmux[1][21] , \outmux[1][20] , \outmux[1][19] , 
        \outmux[1][18] , \outmux[1][17] , \outmux[1][16] , \outmux[1][15] , 
        \outmux[1][14] , \outmux[1][13] , \outmux[1][12] , \outmux[1][11] , 
        \outmux[1][10] , \outmux[1][9] , \outmux[1][8] , \outmux[1][7] , 
        \outmux[1][6] , \outmux[1][5] , \outmux[1][4] , \outmux[1][3] , 
        \outmux[1][2] , \outmux[1][1] , \outmux[1][0] }) );
  mux21N_N32_2 row1_2 ( .in1(in3), .in0(in2), .S(sel[0]), .U({\outmux[2][31] , 
        \outmux[2][30] , \outmux[2][29] , \outmux[2][28] , \outmux[2][27] , 
        \outmux[2][26] , \outmux[2][25] , \outmux[2][24] , \outmux[2][23] , 
        \outmux[2][22] , \outmux[2][21] , \outmux[2][20] , \outmux[2][19] , 
        \outmux[2][18] , \outmux[2][17] , \outmux[2][16] , \outmux[2][15] , 
        \outmux[2][14] , \outmux[2][13] , \outmux[2][12] , \outmux[2][11] , 
        \outmux[2][10] , \outmux[2][9] , \outmux[2][8] , \outmux[2][7] , 
        \outmux[2][6] , \outmux[2][5] , \outmux[2][4] , \outmux[2][3] , 
        \outmux[2][2] , \outmux[2][1] , \outmux[2][0] }) );
  mux21N_N32_1 row2_1 ( .in1({\outmux[2][31] , \outmux[2][30] , 
        \outmux[2][29] , \outmux[2][28] , \outmux[2][27] , \outmux[2][26] , 
        \outmux[2][25] , \outmux[2][24] , \outmux[2][23] , \outmux[2][22] , 
        \outmux[2][21] , \outmux[2][20] , \outmux[2][19] , \outmux[2][18] , 
        \outmux[2][17] , \outmux[2][16] , \outmux[2][15] , \outmux[2][14] , 
        \outmux[2][13] , \outmux[2][12] , \outmux[2][11] , \outmux[2][10] , 
        \outmux[2][9] , \outmux[2][8] , \outmux[2][7] , \outmux[2][6] , 
        \outmux[2][5] , \outmux[2][4] , \outmux[2][3] , \outmux[2][2] , 
        \outmux[2][1] , \outmux[2][0] }), .in0({\outmux[1][31] , 
        \outmux[1][30] , \outmux[1][29] , \outmux[1][28] , \outmux[1][27] , 
        \outmux[1][26] , \outmux[1][25] , \outmux[1][24] , \outmux[1][23] , 
        \outmux[1][22] , \outmux[1][21] , \outmux[1][20] , \outmux[1][19] , 
        \outmux[1][18] , \outmux[1][17] , \outmux[1][16] , \outmux[1][15] , 
        \outmux[1][14] , \outmux[1][13] , \outmux[1][12] , \outmux[1][11] , 
        \outmux[1][10] , \outmux[1][9] , \outmux[1][8] , \outmux[1][7] , 
        \outmux[1][6] , \outmux[1][5] , \outmux[1][4] , \outmux[1][3] , 
        \outmux[1][2] , \outmux[1][1] , \outmux[1][0] }), .S(sel[1]), .U(Y) );
endmodule


module FD_EN_432 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module RegEn_Nbit5_1 ( A, Clk, Reset, EN, U );
  input [4:0] A;
  output [4:0] U;
  input Clk, Reset, EN;


  FD_EN_5 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_4 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_3 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_2 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_1 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
endmodule


module mux21N_N32_7 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   n21, n22, n23, n24;
  assign n21 = S;

  MUX21_399 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n22), .Y(U[0]) );
  MUX21_398 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n22), .Y(U[1]) );
  MUX21_397 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n22), .Y(U[2]) );
  MUX21_396 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n22), .Y(U[3]) );
  MUX21_395 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n22), .Y(U[4]) );
  MUX21_394 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n22), .Y(U[5]) );
  MUX21_393 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n22), .Y(U[6]) );
  MUX21_392 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n22), .Y(U[7]) );
  MUX21_391 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n22), .Y(U[8]) );
  MUX21_390 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n22), .Y(U[9]) );
  MUX21_389 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n22), .Y(U[10]) );
  MUX21_388 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n22), .Y(U[11]) );
  MUX21_387 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n23), .Y(U[12]) );
  MUX21_386 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n23), .Y(U[13]) );
  MUX21_385 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n23), .Y(U[14]) );
  MUX21_384 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n23), .Y(U[15]) );
  MUX21_383 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n23), .Y(U[16]) );
  MUX21_382 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n23), .Y(U[17]) );
  MUX21_381 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n23), .Y(U[18]) );
  MUX21_380 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n23), .Y(U[19]) );
  MUX21_379 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n23), .Y(U[20]) );
  MUX21_378 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n23), .Y(U[21]) );
  MUX21_377 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n23), .Y(U[22]) );
  MUX21_376 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n23), .Y(U[23]) );
  MUX21_375 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n24), .Y(U[24]) );
  MUX21_374 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n24), .Y(U[25]) );
  MUX21_373 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n24), .Y(U[26]) );
  MUX21_372 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n24), .Y(U[27]) );
  MUX21_371 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n24), .Y(U[28]) );
  MUX21_370 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n24), .Y(U[29]) );
  MUX21_369 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n24), .Y(U[30]) );
  MUX21_368 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n24), .Y(U[31]) );
  BUF_X1 U1 ( .A(n21), .Z(n22) );
  BUF_X1 U2 ( .A(n21), .Z(n23) );
  BUF_X1 U3 ( .A(n21), .Z(n24) );
endmodule


module mux21N_N32_8 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   n21, n22, n23, n24;
  assign n21 = S;

  MUX21_431 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n22), .Y(U[0]) );
  MUX21_430 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n22), .Y(U[1]) );
  MUX21_429 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n22), .Y(U[2]) );
  MUX21_428 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n22), .Y(U[3]) );
  MUX21_427 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n22), .Y(U[4]) );
  MUX21_426 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n22), .Y(U[5]) );
  MUX21_425 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n22), .Y(U[6]) );
  MUX21_424 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n22), .Y(U[7]) );
  MUX21_423 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n22), .Y(U[8]) );
  MUX21_422 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n22), .Y(U[9]) );
  MUX21_421 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n22), .Y(U[10]) );
  MUX21_420 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n22), .Y(U[11]) );
  MUX21_419 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n23), .Y(U[12]) );
  MUX21_418 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n23), .Y(U[13]) );
  MUX21_417 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n23), .Y(U[14]) );
  MUX21_416 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n23), .Y(U[15]) );
  MUX21_415 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n23), .Y(U[16]) );
  MUX21_414 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n23), .Y(U[17]) );
  MUX21_413 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n23), .Y(U[18]) );
  MUX21_412 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n23), .Y(U[19]) );
  MUX21_411 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n23), .Y(U[20]) );
  MUX21_410 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n23), .Y(U[21]) );
  MUX21_409 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n23), .Y(U[22]) );
  MUX21_408 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n23), .Y(U[23]) );
  MUX21_407 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n24), .Y(U[24]) );
  MUX21_406 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n24), .Y(U[25]) );
  MUX21_405 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n24), .Y(U[26]) );
  MUX21_404 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n24), .Y(U[27]) );
  MUX21_403 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n24), .Y(U[28]) );
  MUX21_402 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n24), .Y(U[29]) );
  MUX21_401 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n24), .Y(U[30]) );
  MUX21_400 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n24), .Y(U[31]) );
  BUF_X1 U1 ( .A(n21), .Z(n22) );
  BUF_X1 U2 ( .A(n21), .Z(n23) );
  BUF_X1 U3 ( .A(n21), .Z(n24) );
endmodule


module FD_EN_433 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  INV_X1 U3 ( .A(EN), .ZN(n3) );
  NOR2_X1 U4 ( .A1(n2), .A2(RESET), .ZN(n4) );
  AOI22_X1 U5 ( .A1(D), .A2(EN), .B1(n3), .B2(Q), .ZN(n2) );
endmodule


module RegEn_Nbit5_2 ( A, Clk, Reset, EN, U );
  input [4:0] A;
  output [4:0] U;
  input Clk, Reset, EN;


  FD_EN_74 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_73 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_72 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_71 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_70 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
endmodule


module RegEn_Nbit32_3 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;


  FD_EN_106 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_105 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_104 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_103 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_102 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
  FD_EN_101 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[5]) );
  FD_EN_100 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[6]) );
  FD_EN_99 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[7]) );
  FD_EN_98 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[8]) );
  FD_EN_97 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[9]) );
  FD_EN_96 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[10]) );
  FD_EN_95 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[11]) );
  FD_EN_94 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[12]) );
  FD_EN_93 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[13]) );
  FD_EN_92 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[14]) );
  FD_EN_91 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[15]) );
  FD_EN_90 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[16]) );
  FD_EN_89 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[17]) );
  FD_EN_88 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[18]) );
  FD_EN_87 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[19]) );
  FD_EN_86 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[20]) );
  FD_EN_85 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[21]) );
  FD_EN_84 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[22]) );
  FD_EN_83 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[23]) );
  FD_EN_82 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[24]) );
  FD_EN_81 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[25]) );
  FD_EN_80 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[26]) );
  FD_EN_79 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[27]) );
  FD_EN_78 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[28]) );
  FD_EN_77 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[29]) );
  FD_EN_76 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[30]) );
  FD_EN_75 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[31]) );
endmodule


module RegEn_Nbit32_4 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;


  FD_EN_138 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_137 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_136 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_135 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_134 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
  FD_EN_133 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[5]) );
  FD_EN_132 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[6]) );
  FD_EN_131 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[7]) );
  FD_EN_130 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[8]) );
  FD_EN_129 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[9]) );
  FD_EN_128 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[10])
         );
  FD_EN_127 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[11])
         );
  FD_EN_126 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[12])
         );
  FD_EN_125 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[13])
         );
  FD_EN_124 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[14])
         );
  FD_EN_123 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[15])
         );
  FD_EN_122 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[16])
         );
  FD_EN_121 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[17])
         );
  FD_EN_120 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[18])
         );
  FD_EN_119 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[19])
         );
  FD_EN_118 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[20])
         );
  FD_EN_117 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[21])
         );
  FD_EN_116 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[22])
         );
  FD_EN_115 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[23])
         );
  FD_EN_114 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[24])
         );
  FD_EN_113 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[25])
         );
  FD_EN_112 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[26])
         );
  FD_EN_111 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[27])
         );
  FD_EN_110 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[28])
         );
  FD_EN_109 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[29])
         );
  FD_EN_108 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[30])
         );
  FD_EN_107 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[31])
         );
endmodule


module FD_EN_434 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n6, n2, n3;

  DFF_X1 Q_reg ( .D(n6), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n2), .ZN(n6) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module mux81 ( in7, in6, in5, in4, in3, in2, in1, in0, sel, Y );
  input [2:0] sel;
  input in7, in6, in5, in4, in3, in2, in1, in0;
  output Y;

  wire   [4:1] outmux;
  wire   [2:1] outmux2;
  tri   [2:0] sel;

  MUX21_438 row1_1 ( .in1(in1), .in0(in0), .S(sel[0]), .Y(outmux[1]) );
  MUX21_437 row1_2 ( .in1(in3), .in0(in2), .S(sel[0]), .Y(outmux[2]) );
  MUX21_436 row1_3 ( .in1(in5), .in0(in4), .S(sel[0]), .Y(outmux[3]) );
  MUX21_435 row1_4 ( .in1(in7), .in0(in6), .S(sel[0]), .Y(outmux[4]) );
  MUX21_434 row2_1 ( .in1(outmux[2]), .in0(outmux[1]), .S(sel[1]), .Y(
        outmux2[1]) );
  MUX21_433 row2_2 ( .in1(outmux[4]), .in0(outmux[3]), .S(sel[1]), .Y(
        outmux2[2]) );
  MUX21_432 row3_1 ( .in1(outmux2[2]), .in0(outmux2[1]), .S(sel[2]), .Y(Y) );
endmodule


module ALU_v2 ( A, B, ALUsel, unsign, arith_logN, ALUout, AeqB, AnoteqB, AgB, 
        AlB, AgeqB, AleqB );
  input [31:0] A;
  input [31:0] B;
  input [3:0] ALUsel;
  output [31:0] ALUout;
  input unsign, arith_logN;
  output AeqB, AnoteqB, AgB, AlB, AgeqB, AleqB;
  wire   AinMUL_0_port, AinMUL_1_port, AinMUL_2_port, AinMUL_3_port,
         AinMUL_4_port, AinMUL_5_port, AinMUL_6_port, AinMUL_7_port,
         AinMUL_8_port, AinMUL_9_port, AinMUL_10_port, AinMUL_11_port,
         AinMUL_12_port, AinMUL_13_port, AinMUL_14_port, AinMUL_15_port,
         BinMUL_0_port, BinMUL_1_port, BinMUL_2_port, BinMUL_3_port,
         BinMUL_4_port, BinMUL_5_port, BinMUL_6_port, BinMUL_7_port,
         BinMUL_8_port, BinMUL_9_port, BinMUL_10_port, BinMUL_11_port,
         BinMUL_12_port, BinMUL_13_port, BinMUL_14_port, BinMUL_15_port,
         MULout_0_port, MULout_1_port, MULout_2_port, MULout_3_port,
         MULout_4_port, MULout_5_port, MULout_6_port, MULout_7_port,
         MULout_8_port, MULout_9_port, MULout_10_port, MULout_11_port,
         MULout_12_port, MULout_13_port, MULout_14_port, MULout_15_port,
         MULout_16_port, MULout_17_port, MULout_18_port, MULout_19_port,
         MULout_20_port, MULout_21_port, MULout_22_port, MULout_23_port,
         MULout_24_port, MULout_25_port, MULout_26_port, MULout_27_port,
         MULout_28_port, MULout_29_port, MULout_30_port, MULout_31_port,
         AinADDSUB_0_port, AinADDSUB_1_port, AinADDSUB_2_port,
         AinADDSUB_3_port, AinADDSUB_4_port, AinADDSUB_5_port,
         AinADDSUB_6_port, AinADDSUB_7_port, AinADDSUB_8_port,
         AinADDSUB_9_port, AinADDSUB_10_port, AinADDSUB_11_port,
         AinADDSUB_12_port, AinADDSUB_13_port, AinADDSUB_14_port,
         AinADDSUB_15_port, AinADDSUB_16_port, AinADDSUB_17_port,
         AinADDSUB_18_port, AinADDSUB_19_port, AinADDSUB_20_port,
         AinADDSUB_21_port, AinADDSUB_22_port, AinADDSUB_23_port,
         AinADDSUB_24_port, AinADDSUB_25_port, AinADDSUB_26_port,
         AinADDSUB_27_port, AinADDSUB_28_port, AinADDSUB_29_port,
         AinADDSUB_30_port, AinADDSUB_31_port, BinADDSUB_0_port,
         BinADDSUB_1_port, BinADDSUB_2_port, BinADDSUB_3_port,
         BinADDSUB_4_port, BinADDSUB_5_port, BinADDSUB_6_port,
         BinADDSUB_7_port, BinADDSUB_8_port, BinADDSUB_9_port,
         BinADDSUB_10_port, BinADDSUB_11_port, BinADDSUB_12_port,
         BinADDSUB_13_port, BinADDSUB_14_port, BinADDSUB_15_port,
         BinADDSUB_16_port, BinADDSUB_17_port, BinADDSUB_18_port,
         BinADDSUB_19_port, BinADDSUB_20_port, BinADDSUB_21_port,
         BinADDSUB_22_port, BinADDSUB_23_port, BinADDSUB_24_port,
         BinADDSUB_25_port, BinADDSUB_26_port, BinADDSUB_27_port,
         BinADDSUB_28_port, BinADDSUB_29_port, BinADDSUB_30_port,
         BinADDSUB_31_port, ADDSUBout_0_port, ADDSUBout_1_port,
         ADDSUBout_2_port, ADDSUBout_3_port, ADDSUBout_4_port,
         ADDSUBout_5_port, ADDSUBout_6_port, ADDSUBout_7_port,
         ADDSUBout_8_port, ADDSUBout_9_port, ADDSUBout_10_port,
         ADDSUBout_11_port, ADDSUBout_12_port, ADDSUBout_13_port,
         ADDSUBout_14_port, ADDSUBout_15_port, ADDSUBout_16_port,
         ADDSUBout_17_port, ADDSUBout_18_port, ADDSUBout_19_port,
         ADDSUBout_20_port, ADDSUBout_21_port, ADDSUBout_22_port,
         ADDSUBout_23_port, ADDSUBout_24_port, ADDSUBout_25_port,
         ADDSUBout_26_port, ADDSUBout_27_port, ADDSUBout_28_port,
         ADDSUBout_29_port, ADDSUBout_30_port, ADDSUBout_31_port, sumnsub,
         Carry, AinLOGIC_0_port, AinLOGIC_1_port, AinLOGIC_2_port,
         AinLOGIC_3_port, AinLOGIC_4_port, AinLOGIC_5_port, AinLOGIC_6_port,
         AinLOGIC_7_port, AinLOGIC_8_port, AinLOGIC_9_port, AinLOGIC_10_port,
         AinLOGIC_11_port, AinLOGIC_12_port, AinLOGIC_13_port,
         AinLOGIC_14_port, AinLOGIC_15_port, AinLOGIC_16_port,
         AinLOGIC_17_port, AinLOGIC_18_port, AinLOGIC_19_port,
         AinLOGIC_20_port, AinLOGIC_21_port, AinLOGIC_22_port,
         AinLOGIC_23_port, AinLOGIC_24_port, AinLOGIC_25_port,
         AinLOGIC_26_port, AinLOGIC_27_port, AinLOGIC_28_port,
         AinLOGIC_29_port, AinLOGIC_30_port, AinLOGIC_31_port, BinLOGIC_0_port,
         BinLOGIC_1_port, BinLOGIC_2_port, BinLOGIC_3_port, BinLOGIC_4_port,
         BinLOGIC_5_port, BinLOGIC_6_port, BinLOGIC_7_port, BinLOGIC_8_port,
         BinLOGIC_9_port, BinLOGIC_10_port, BinLOGIC_11_port, BinLOGIC_12_port,
         BinLOGIC_13_port, BinLOGIC_14_port, BinLOGIC_15_port,
         BinLOGIC_16_port, BinLOGIC_17_port, BinLOGIC_18_port,
         BinLOGIC_19_port, BinLOGIC_20_port, BinLOGIC_21_port,
         BinLOGIC_22_port, BinLOGIC_23_port, BinLOGIC_24_port,
         BinLOGIC_25_port, BinLOGIC_26_port, BinLOGIC_27_port,
         BinLOGIC_28_port, BinLOGIC_29_port, BinLOGIC_30_port,
         BinLOGIC_31_port, notAout_0_port, notAout_1_port, notAout_2_port,
         notAout_3_port, notAout_4_port, notAout_5_port, notAout_6_port,
         notAout_7_port, notAout_8_port, notAout_9_port, notAout_10_port,
         notAout_11_port, notAout_12_port, notAout_13_port, notAout_14_port,
         notAout_15_port, notAout_16_port, notAout_17_port, notAout_18_port,
         notAout_19_port, notAout_20_port, notAout_21_port, notAout_22_port,
         notAout_23_port, notAout_24_port, notAout_25_port, notAout_26_port,
         notAout_27_port, notAout_28_port, notAout_29_port, notAout_30_port,
         notAout_31_port, notBout_0_port, notBout_1_port, notBout_2_port,
         notBout_3_port, notBout_4_port, notBout_5_port, notBout_6_port,
         notBout_7_port, notBout_8_port, notBout_9_port, notBout_10_port,
         notBout_11_port, notBout_12_port, notBout_13_port, notBout_14_port,
         notBout_15_port, notBout_16_port, notBout_17_port, notBout_18_port,
         notBout_19_port, notBout_20_port, notBout_21_port, notBout_22_port,
         notBout_23_port, notBout_24_port, notBout_25_port, notBout_26_port,
         notBout_27_port, notBout_28_port, notBout_29_port, notBout_30_port,
         notBout_31_port, AorBout_0_port, AorBout_1_port, AorBout_2_port,
         AorBout_3_port, AorBout_4_port, AorBout_5_port, AorBout_6_port,
         AorBout_7_port, AorBout_8_port, AorBout_9_port, AorBout_10_port,
         AorBout_11_port, AorBout_12_port, AorBout_13_port, AorBout_14_port,
         AorBout_15_port, AorBout_16_port, AorBout_17_port, AorBout_18_port,
         AorBout_19_port, AorBout_20_port, AorBout_21_port, AorBout_22_port,
         AorBout_23_port, AorBout_24_port, AorBout_25_port, AorBout_26_port,
         AorBout_27_port, AorBout_28_port, AorBout_29_port, AorBout_30_port,
         AorBout_31_port, AxorBout_0_port, AxorBout_1_port, AxorBout_2_port,
         AxorBout_3_port, AxorBout_4_port, AxorBout_5_port, AxorBout_6_port,
         AxorBout_7_port, AxorBout_8_port, AxorBout_9_port, AxorBout_10_port,
         AxorBout_11_port, AxorBout_12_port, AxorBout_13_port,
         AxorBout_14_port, AxorBout_15_port, AxorBout_16_port,
         AxorBout_17_port, AxorBout_18_port, AxorBout_19_port,
         AxorBout_20_port, AxorBout_21_port, AxorBout_22_port,
         AxorBout_23_port, AxorBout_24_port, AxorBout_25_port,
         AxorBout_26_port, AxorBout_27_port, AxorBout_28_port,
         AxorBout_29_port, AxorBout_30_port, AxorBout_31_port, N1020, N1021,
         Right_LeftN, N1008, N1009, enADDSUB, enMUL, N1015, enLOGIC, N1017,
         enSHIFTER, N1019, Shift_Rotaten, N945, N947, N949, N951, N953, N955,
         N957, N959, N961, N963, N965, N967, N969, N971, N973, N975, N977,
         N979, N981, N983, N985, N987, N989, N991, N993, N995, N997, N999,
         N1001, N1003, N1005, N1007, AinSHIFTER_0_port, AinSHIFTER_1_port,
         AinSHIFTER_2_port, AinSHIFTER_3_port, AinSHIFTER_4_port,
         AinSHIFTER_5_port, AinSHIFTER_6_port, AinSHIFTER_7_port,
         AinSHIFTER_8_port, AinSHIFTER_9_port, AinSHIFTER_10_port,
         AinSHIFTER_11_port, AinSHIFTER_12_port, AinSHIFTER_13_port,
         AinSHIFTER_14_port, AinSHIFTER_15_port, AinSHIFTER_16_port,
         AinSHIFTER_17_port, AinSHIFTER_18_port, AinSHIFTER_19_port,
         AinSHIFTER_20_port, AinSHIFTER_21_port, AinSHIFTER_22_port,
         AinSHIFTER_23_port, AinSHIFTER_24_port, AinSHIFTER_25_port,
         AinSHIFTER_26_port, AinSHIFTER_27_port, AinSHIFTER_28_port,
         AinSHIFTER_29_port, AinSHIFTER_30_port, AinSHIFTER_31_port,
         Binshift_0_port, Binshift_1_port, Binshift_2_port, Binshift_3_port,
         Binshift_4_port, SHIFTERout_0_port, SHIFTERout_1_port,
         SHIFTERout_2_port, SHIFTERout_3_port, SHIFTERout_4_port,
         SHIFTERout_5_port, SHIFTERout_6_port, SHIFTERout_7_port,
         SHIFTERout_8_port, SHIFTERout_9_port, SHIFTERout_10_port,
         SHIFTERout_11_port, SHIFTERout_12_port, SHIFTERout_13_port,
         SHIFTERout_14_port, SHIFTERout_15_port, SHIFTERout_16_port,
         SHIFTERout_17_port, SHIFTERout_18_port, SHIFTERout_19_port,
         SHIFTERout_20_port, SHIFTERout_21_port, SHIFTERout_22_port,
         SHIFTERout_23_port, SHIFTERout_24_port, SHIFTERout_25_port,
         SHIFTERout_26_port, SHIFTERout_27_port, SHIFTERout_28_port,
         SHIFTERout_29_port, SHIFTERout_30_port, SHIFTERout_31_port, complete,
         n336, n342, n345, n352, n355, n361, n364, n370, n373, n379, n382,
         n388, n391, n397, n400, n406, n409, n421, n424, n430, n433, n439,
         n442, n448, n451, n452, n454, n455, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n1069, n1072,
         n1076, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n92, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n324, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n337, n338, n339, n340, n341, n343,
         n344, n346, n347, n348, n349, n350, n351, n353, n354, n356, n357,
         n358, n359, n360, n362, n363, n365, n366, n367, n368, n369, n371,
         n372, n374, n375, n376, n377, n378, n380, n381, n383, n384, n385,
         n386, n387, n389, n390, n392, n393, n394, n395, n396, n398, n399,
         n401, n402, n403, n404, n405, n407, n408, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n422, n423, n425, n426,
         n427, n428, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136;
  tri   [3:0] ALUsel;
  tri   unsign;
  tri   arith_logN;

  DLH_X1 Right_LeftN_reg ( .G(N1020), .D(N1021), .Q(Right_LeftN) );
  DLH_X1 enADDSUB_reg ( .G(n1127), .D(n1133), .Q(enADDSUB) );
  DLH_X1 enMUL_reg ( .G(n1127), .D(n1136), .Q(enMUL) );
  DLH_X1 enLOGIC_reg ( .G(n1127), .D(N1015), .Q(enLOGIC) );
  DLH_X1 enSHIFTER_reg ( .G(n1127), .D(N1017), .Q(enSHIFTER) );
  DLH_X1 Shift_Rotaten_reg ( .G(n1130), .D(N1019), .Q(Shift_Rotaten) );
  DLH_X1 ALUout_reg_0_inst ( .G(n1128), .D(N945), .Q(ALUout[0]) );
  DLH_X1 ALUout_reg_1_inst ( .G(n1127), .D(N947), .Q(ALUout[1]) );
  DLH_X1 ALUout_reg_2_inst ( .G(n1127), .D(N949), .Q(ALUout[2]) );
  DLH_X1 ALUout_reg_3_inst ( .G(n1130), .D(N951), .Q(ALUout[3]) );
  DLH_X1 ALUout_reg_4_inst ( .G(n1129), .D(N953), .Q(ALUout[4]) );
  DLH_X1 ALUout_reg_5_inst ( .G(n1130), .D(N955), .Q(ALUout[5]) );
  DLH_X1 ALUout_reg_6_inst ( .G(n1129), .D(N957), .Q(ALUout[6]) );
  DLH_X1 ALUout_reg_7_inst ( .G(n1129), .D(N959), .Q(ALUout[7]) );
  DLH_X1 ALUout_reg_8_inst ( .G(n1129), .D(N961), .Q(ALUout[8]) );
  DLH_X1 ALUout_reg_9_inst ( .G(n1129), .D(N963), .Q(ALUout[9]) );
  DLH_X1 ALUout_reg_10_inst ( .G(n1127), .D(N965), .Q(ALUout[10]) );
  DLH_X1 ALUout_reg_11_inst ( .G(n1127), .D(N967), .Q(ALUout[11]) );
  DLH_X1 ALUout_reg_12_inst ( .G(n1129), .D(N969), .Q(ALUout[12]) );
  DLH_X1 ALUout_reg_13_inst ( .G(n1129), .D(N971), .Q(ALUout[13]) );
  DLH_X1 ALUout_reg_14_inst ( .G(n1129), .D(N973), .Q(ALUout[14]) );
  DLH_X1 ALUout_reg_15_inst ( .G(n1130), .D(N975), .Q(ALUout[15]) );
  DLH_X1 ALUout_reg_16_inst ( .G(n1128), .D(N977), .Q(ALUout[16]) );
  DLH_X1 ALUout_reg_17_inst ( .G(n1128), .D(N979), .Q(ALUout[17]) );
  DLH_X1 ALUout_reg_18_inst ( .G(n1128), .D(N981), .Q(ALUout[18]) );
  DLH_X1 ALUout_reg_19_inst ( .G(n1128), .D(N983), .Q(ALUout[19]) );
  DLH_X1 ALUout_reg_20_inst ( .G(n1127), .D(N985), .Q(ALUout[20]) );
  DLH_X1 ALUout_reg_21_inst ( .G(n1127), .D(N987), .Q(ALUout[21]) );
  DLH_X1 ALUout_reg_22_inst ( .G(n1128), .D(N989), .Q(ALUout[22]) );
  DLH_X1 ALUout_reg_23_inst ( .G(n1128), .D(N991), .Q(ALUout[23]) );
  DLH_X1 ALUout_reg_24_inst ( .G(n1128), .D(N993), .Q(ALUout[24]) );
  DLH_X1 ALUout_reg_25_inst ( .G(n1128), .D(N995), .Q(ALUout[25]) );
  DLH_X1 ALUout_reg_26_inst ( .G(n1128), .D(N997), .Q(ALUout[26]) );
  DLH_X1 ALUout_reg_27_inst ( .G(n1128), .D(N999), .Q(ALUout[27]) );
  DLH_X1 ALUout_reg_28_inst ( .G(n1127), .D(N1001), .Q(ALUout[28]) );
  DLH_X1 ALUout_reg_29_inst ( .G(n1129), .D(N1003), .Q(ALUout[29]) );
  DLH_X1 ALUout_reg_30_inst ( .G(n1129), .D(N1005), .Q(ALUout[30]) );
  DLH_X1 ALUout_reg_31_inst ( .G(n1129), .D(N1007), .Q(ALUout[31]) );
  BoothMulWallace_Nbit32 MUL ( .a({AinMUL_15_port, AinMUL_14_port, 
        AinMUL_13_port, AinMUL_12_port, AinMUL_11_port, AinMUL_10_port, 
        AinMUL_9_port, AinMUL_8_port, AinMUL_7_port, AinMUL_6_port, 
        AinMUL_5_port, AinMUL_4_port, AinMUL_3_port, AinMUL_2_port, 
        AinMUL_1_port, AinMUL_0_port}), .b({BinMUL_15_port, BinMUL_14_port, 
        BinMUL_13_port, BinMUL_12_port, BinMUL_11_port, BinMUL_10_port, 
        BinMUL_9_port, BinMUL_8_port, BinMUL_7_port, BinMUL_6_port, 
        BinMUL_5_port, BinMUL_4_port, BinMUL_3_port, BinMUL_2_port, 
        BinMUL_1_port, BinMUL_0_port}), .p({MULout_31_port, MULout_30_port, 
        MULout_29_port, MULout_28_port, MULout_27_port, MULout_26_port, 
        MULout_25_port, MULout_24_port, MULout_23_port, MULout_22_port, 
        MULout_21_port, MULout_20_port, MULout_19_port, MULout_18_port, 
        MULout_17_port, MULout_16_port, MULout_15_port, MULout_14_port, 
        MULout_13_port, MULout_12_port, MULout_11_port, MULout_10_port, 
        MULout_9_port, MULout_8_port, MULout_7_port, MULout_6_port, 
        MULout_5_port, MULout_4_port, MULout_3_port, MULout_2_port, 
        MULout_1_port, MULout_0_port}) );
  AddSubN_Nbit32_1 ADDSUB ( .A({AinADDSUB_31_port, AinADDSUB_30_port, 
        AinADDSUB_29_port, AinADDSUB_28_port, AinADDSUB_27_port, 
        AinADDSUB_26_port, AinADDSUB_25_port, AinADDSUB_24_port, 
        AinADDSUB_23_port, AinADDSUB_22_port, AinADDSUB_21_port, 
        AinADDSUB_20_port, AinADDSUB_19_port, AinADDSUB_18_port, 
        AinADDSUB_17_port, AinADDSUB_16_port, AinADDSUB_15_port, 
        AinADDSUB_14_port, AinADDSUB_13_port, AinADDSUB_12_port, 
        AinADDSUB_11_port, AinADDSUB_10_port, AinADDSUB_9_port, 
        AinADDSUB_8_port, AinADDSUB_7_port, AinADDSUB_6_port, AinADDSUB_5_port, 
        AinADDSUB_4_port, AinADDSUB_3_port, AinADDSUB_2_port, AinADDSUB_1_port, 
        AinADDSUB_0_port}), .B({BinADDSUB_31_port, BinADDSUB_30_port, 
        BinADDSUB_29_port, BinADDSUB_28_port, BinADDSUB_27_port, 
        BinADDSUB_26_port, BinADDSUB_25_port, BinADDSUB_24_port, 
        BinADDSUB_23_port, BinADDSUB_22_port, BinADDSUB_21_port, 
        BinADDSUB_20_port, BinADDSUB_19_port, BinADDSUB_18_port, 
        BinADDSUB_17_port, BinADDSUB_16_port, BinADDSUB_15_port, 
        BinADDSUB_14_port, BinADDSUB_13_port, BinADDSUB_12_port, 
        BinADDSUB_11_port, BinADDSUB_10_port, BinADDSUB_9_port, 
        BinADDSUB_8_port, BinADDSUB_7_port, BinADDSUB_6_port, BinADDSUB_5_port, 
        BinADDSUB_4_port, BinADDSUB_3_port, BinADDSUB_2_port, BinADDSUB_1_port, 
        BinADDSUB_0_port}), .addnsub(sumnsub), .S({ADDSUBout_31_port, 
        ADDSUBout_30_port, ADDSUBout_29_port, ADDSUBout_28_port, 
        ADDSUBout_27_port, ADDSUBout_26_port, ADDSUBout_25_port, 
        ADDSUBout_24_port, ADDSUBout_23_port, ADDSUBout_22_port, 
        ADDSUBout_21_port, ADDSUBout_20_port, ADDSUBout_19_port, 
        ADDSUBout_18_port, ADDSUBout_17_port, ADDSUBout_16_port, 
        ADDSUBout_15_port, ADDSUBout_14_port, ADDSUBout_13_port, 
        ADDSUBout_12_port, ADDSUBout_11_port, ADDSUBout_10_port, 
        ADDSUBout_9_port, ADDSUBout_8_port, ADDSUBout_7_port, ADDSUBout_6_port, 
        ADDSUBout_5_port, ADDSUBout_4_port, ADDSUBout_3_port, ADDSUBout_2_port, 
        ADDSUBout_1_port, ADDSUBout_0_port}), .Cout(Carry) );
  Comp_Nbit32 COMPLog ( .signA(AinADDSUB_31_port), .signB(BinADDSUB_31_port), 
        .Diff({ADDSUBout_31_port, ADDSUBout_30_port, ADDSUBout_29_port, 
        ADDSUBout_28_port, ADDSUBout_27_port, ADDSUBout_26_port, 
        ADDSUBout_25_port, ADDSUBout_24_port, ADDSUBout_23_port, 
        ADDSUBout_22_port, ADDSUBout_21_port, ADDSUBout_20_port, 
        ADDSUBout_19_port, ADDSUBout_18_port, ADDSUBout_17_port, 
        ADDSUBout_16_port, ADDSUBout_15_port, ADDSUBout_14_port, 
        ADDSUBout_13_port, ADDSUBout_12_port, ADDSUBout_11_port, 
        ADDSUBout_10_port, ADDSUBout_9_port, ADDSUBout_8_port, 
        ADDSUBout_7_port, ADDSUBout_6_port, ADDSUBout_5_port, ADDSUBout_4_port, 
        ADDSUBout_3_port, ADDSUBout_2_port, ADDSUBout_1_port, ADDSUBout_0_port}), .Carry(Carry), .unsign(unsign), .AgB(AgB), .AeqB(AeqB), .AnoteqB(AnoteqB), 
        .AlB(AlB), .AgeqB(AgeqB), .AleqB(AleqB) );
  LogicFun_v2_Nbit32 LOGICunit ( .A({AinLOGIC_31_port, AinLOGIC_30_port, 
        AinLOGIC_29_port, AinLOGIC_28_port, AinLOGIC_27_port, AinLOGIC_26_port, 
        AinLOGIC_25_port, AinLOGIC_24_port, AinLOGIC_23_port, AinLOGIC_22_port, 
        AinLOGIC_21_port, AinLOGIC_20_port, AinLOGIC_19_port, AinLOGIC_18_port, 
        AinLOGIC_17_port, AinLOGIC_16_port, AinLOGIC_15_port, AinLOGIC_14_port, 
        AinLOGIC_13_port, AinLOGIC_12_port, AinLOGIC_11_port, AinLOGIC_10_port, 
        AinLOGIC_9_port, AinLOGIC_8_port, AinLOGIC_7_port, AinLOGIC_6_port, 
        AinLOGIC_5_port, AinLOGIC_4_port, AinLOGIC_3_port, AinLOGIC_2_port, 
        AinLOGIC_1_port, AinLOGIC_0_port}), .B({BinLOGIC_31_port, 
        BinLOGIC_30_port, BinLOGIC_29_port, BinLOGIC_28_port, BinLOGIC_27_port, 
        BinLOGIC_26_port, BinLOGIC_25_port, BinLOGIC_24_port, BinLOGIC_23_port, 
        BinLOGIC_22_port, BinLOGIC_21_port, BinLOGIC_20_port, BinLOGIC_19_port, 
        BinLOGIC_18_port, BinLOGIC_17_port, BinLOGIC_16_port, BinLOGIC_15_port, 
        BinLOGIC_14_port, BinLOGIC_13_port, BinLOGIC_12_port, BinLOGIC_11_port, 
        BinLOGIC_10_port, BinLOGIC_9_port, BinLOGIC_8_port, BinLOGIC_7_port, 
        BinLOGIC_6_port, BinLOGIC_5_port, BinLOGIC_4_port, BinLOGIC_3_port, 
        BinLOGIC_2_port, BinLOGIC_1_port, BinLOGIC_0_port}), .notA({
        notAout_31_port, notAout_30_port, notAout_29_port, notAout_28_port, 
        notAout_27_port, notAout_26_port, notAout_25_port, notAout_24_port, 
        notAout_23_port, notAout_22_port, notAout_21_port, notAout_20_port, 
        notAout_19_port, notAout_18_port, notAout_17_port, notAout_16_port, 
        notAout_15_port, notAout_14_port, notAout_13_port, notAout_12_port, 
        notAout_11_port, notAout_10_port, notAout_9_port, notAout_8_port, 
        notAout_7_port, notAout_6_port, notAout_5_port, notAout_4_port, 
        notAout_3_port, notAout_2_port, notAout_1_port, notAout_0_port}), 
        .notB({notBout_31_port, notBout_30_port, notBout_29_port, 
        notBout_28_port, notBout_27_port, notBout_26_port, notBout_25_port, 
        notBout_24_port, notBout_23_port, notBout_22_port, notBout_21_port, 
        notBout_20_port, notBout_19_port, notBout_18_port, notBout_17_port, 
        notBout_16_port, notBout_15_port, notBout_14_port, notBout_13_port, 
        notBout_12_port, notBout_11_port, notBout_10_port, notBout_9_port, 
        notBout_8_port, notBout_7_port, notBout_6_port, notBout_5_port, 
        notBout_4_port, notBout_3_port, notBout_2_port, notBout_1_port, 
        notBout_0_port}), .AandB({n345, n388, n391, n352, n364, n370, n373, 
        n336, n379, n382, n342, n355, n361, n406, n409, n421, n424, n430, n539, 
        n540, n538, n541, n433, n439, n442, n448, n451, n452, n454, n397, n400, 
        n455}), .AorB({AorBout_31_port, AorBout_30_port, AorBout_29_port, 
        AorBout_28_port, AorBout_27_port, AorBout_26_port, AorBout_25_port, 
        AorBout_24_port, AorBout_23_port, AorBout_22_port, AorBout_21_port, 
        AorBout_20_port, AorBout_19_port, AorBout_18_port, AorBout_17_port, 
        AorBout_16_port, AorBout_15_port, AorBout_14_port, AorBout_13_port, 
        AorBout_12_port, AorBout_11_port, AorBout_10_port, AorBout_9_port, 
        AorBout_8_port, AorBout_7_port, AorBout_6_port, AorBout_5_port, 
        AorBout_4_port, AorBout_3_port, AorBout_2_port, AorBout_1_port, 
        AorBout_0_port}), .AxorB({AxorBout_31_port, AxorBout_30_port, 
        AxorBout_29_port, AxorBout_28_port, AxorBout_27_port, AxorBout_26_port, 
        AxorBout_25_port, AxorBout_24_port, AxorBout_23_port, AxorBout_22_port, 
        AxorBout_21_port, AxorBout_20_port, AxorBout_19_port, AxorBout_18_port, 
        AxorBout_17_port, AxorBout_16_port, AxorBout_15_port, AxorBout_14_port, 
        AxorBout_13_port, AxorBout_12_port, AxorBout_11_port, AxorBout_10_port, 
        AxorBout_9_port, AxorBout_8_port, AxorBout_7_port, AxorBout_6_port, 
        AxorBout_5_port, AxorBout_4_port, AxorBout_3_port, AxorBout_2_port, 
        AxorBout_1_port, AxorBout_0_port}), .AnorB({n568, n572, n573, n569, 
        n570, n561, n571, n558, n562, n563, n567, n559, n560, n564, n565, n566, 
        n549, n543, n550, n544, n546, n545, n551, n552, n553, n554, n555, n556, 
        n557, n547, n542, n548}) );
  bidir_shift_rot_N_interface_NBIT32 SHIFTER ( .data_in({AinSHIFTER_31_port, 
        AinSHIFTER_30_port, AinSHIFTER_29_port, AinSHIFTER_28_port, 
        AinSHIFTER_27_port, AinSHIFTER_26_port, AinSHIFTER_25_port, 
        AinSHIFTER_24_port, AinSHIFTER_23_port, AinSHIFTER_22_port, 
        AinSHIFTER_21_port, AinSHIFTER_20_port, AinSHIFTER_19_port, 
        AinSHIFTER_18_port, AinSHIFTER_17_port, AinSHIFTER_16_port, 
        AinSHIFTER_15_port, AinSHIFTER_14_port, AinSHIFTER_13_port, 
        AinSHIFTER_12_port, AinSHIFTER_11_port, AinSHIFTER_10_port, 
        AinSHIFTER_9_port, AinSHIFTER_8_port, AinSHIFTER_7_port, 
        AinSHIFTER_6_port, AinSHIFTER_5_port, AinSHIFTER_4_port, 
        AinSHIFTER_3_port, AinSHIFTER_2_port, AinSHIFTER_1_port, 
        AinSHIFTER_0_port}), .moves({Binshift_4_port, Binshift_3_port, 
        Binshift_2_port, Binshift_1_port, Binshift_0_port}), .tot(complete), 
        .shift_rotN(Shift_Rotaten), .right_leftN(Right_LeftN), .arith_logN(
        arith_logN), .data_out({SHIFTERout_31_port, SHIFTERout_30_port, 
        SHIFTERout_29_port, SHIFTERout_28_port, SHIFTERout_27_port, 
        SHIFTERout_26_port, SHIFTERout_25_port, SHIFTERout_24_port, 
        SHIFTERout_23_port, SHIFTERout_22_port, SHIFTERout_21_port, 
        SHIFTERout_20_port, SHIFTERout_19_port, SHIFTERout_18_port, 
        SHIFTERout_17_port, SHIFTERout_16_port, SHIFTERout_15_port, 
        SHIFTERout_14_port, SHIFTERout_13_port, SHIFTERout_12_port, 
        SHIFTERout_11_port, SHIFTERout_10_port, SHIFTERout_9_port, 
        SHIFTERout_8_port, SHIFTERout_7_port, SHIFTERout_6_port, 
        SHIFTERout_5_port, SHIFTERout_4_port, SHIFTERout_3_port, 
        SHIFTERout_2_port, SHIFTERout_1_port, SHIFTERout_0_port}) );
  DLH_X1 sumnsub_reg ( .G(N1008), .D(N1009), .Q(sumnsub) );
  NAND3_X1 U563 ( .A1(n289), .A2(n290), .A3(N1017), .ZN(N1020) );
  NAND3_X1 U565 ( .A1(n328), .A2(n329), .A3(n81), .ZN(n98) );
  NAND3_X1 U566 ( .A1(ALUsel[1]), .A2(n329), .A3(n81), .ZN(n99) );
  NAND3_X1 U567 ( .A1(n329), .A2(n330), .A3(n328), .ZN(n292) );
  NAND3_X1 U568 ( .A1(n354), .A2(n356), .A3(n357), .ZN(n353) );
  NAND3_X1 U569 ( .A1(n366), .A2(n367), .A3(n368), .ZN(n365) );
  NOR2_X1 U1 ( .A1(n1090), .A2(n427), .ZN(AinADDSUB_10_port) );
  NOR2_X1 U2 ( .A1(n1088), .A2(n402), .ZN(AinADDSUB_2_port) );
  NOR2_X1 U3 ( .A1(n1088), .A2(n398), .ZN(AinADDSUB_3_port) );
  NOR2_X1 U4 ( .A1(n1088), .A2(n404), .ZN(AinADDSUB_28_port) );
  NOR2_X1 U5 ( .A1(n1088), .A2(n405), .ZN(AinADDSUB_27_port) );
  INV_X1 U6 ( .A(A[2]), .ZN(n402) );
  INV_X1 U7 ( .A(A[3]), .ZN(n398) );
  INV_X1 U8 ( .A(A[9]), .ZN(n390) );
  INV_X1 U9 ( .A(A[10]), .ZN(n427) );
  INV_X1 U10 ( .A(A[11]), .ZN(n426) );
  INV_X1 U11 ( .A(A[13]), .ZN(n423) );
  INV_X1 U12 ( .A(A[14]), .ZN(n422) );
  INV_X1 U13 ( .A(A[15]), .ZN(n420) );
  BUF_X1 U14 ( .A(n387), .Z(n1087) );
  NOR2_X1 U15 ( .A1(n1087), .A2(n390), .ZN(AinADDSUB_9_port) );
  BUF_X1 U16 ( .A(n85), .Z(n1124) );
  BUF_X1 U17 ( .A(n85), .Z(n1125) );
  BUF_X1 U18 ( .A(n85), .Z(n1126) );
  AND2_X1 U19 ( .A1(n1126), .A2(n1108), .ZN(N1017) );
  NOR3_X1 U20 ( .A1(n1123), .A2(n1136), .A3(n1131), .ZN(n85) );
  BUF_X1 U21 ( .A(n96), .Z(n1106) );
  BUF_X1 U22 ( .A(n96), .Z(n1107) );
  BUF_X1 U23 ( .A(n1072), .Z(n1132) );
  BUF_X1 U24 ( .A(n96), .Z(n1108) );
  BUF_X1 U25 ( .A(n1072), .Z(n1133) );
  BUF_X1 U26 ( .A(n1072), .Z(n1131) );
  AOI221_X1 U27 ( .B1(notBout_25_port), .B2(n1120), .C1(n373), .C2(n1116), .A(
        n112), .ZN(n111) );
  OAI22_X1 U28 ( .A1(AorBout_25_port), .A2(n1114), .B1(n571), .B2(n1113), .ZN(
        n112) );
  AOI221_X1 U29 ( .B1(notBout_31_port), .B2(n1118), .C1(n345), .C2(n1116), .A(
        n300), .ZN(n299) );
  OAI22_X1 U30 ( .A1(AorBout_31_port), .A2(n1114), .B1(n568), .B2(n1112), .ZN(
        n300) );
  AOI221_X1 U31 ( .B1(notBout_29_port), .B2(n1118), .C1(n391), .C2(n1116), .A(
        n314), .ZN(n313) );
  OAI22_X1 U32 ( .A1(AorBout_29_port), .A2(n1114), .B1(n573), .B2(n1113), .ZN(
        n314) );
  AOI221_X1 U33 ( .B1(notBout_28_port), .B2(n1118), .C1(n352), .C2(n1116), .A(
        n321), .ZN(n320) );
  OAI22_X1 U34 ( .A1(AorBout_28_port), .A2(n1114), .B1(n569), .B2(n1112), .ZN(
        n321) );
  NOR2_X1 U35 ( .A1(n1093), .A2(n381), .ZN(BinLOGIC_24_port) );
  NOR2_X1 U36 ( .A1(n1093), .A2(n383), .ZN(BinLOGIC_23_port) );
  NOR2_X1 U37 ( .A1(n1093), .A2(n384), .ZN(BinLOGIC_18_port) );
  NOR2_X1 U38 ( .A1(n1093), .A2(n385), .ZN(BinLOGIC_17_port) );
  NOR2_X1 U39 ( .A1(n1093), .A2(n386), .ZN(BinLOGIC_16_port) );
  NOR2_X1 U40 ( .A1(n1092), .A2(n378), .ZN(BinLOGIC_29_port) );
  NOR2_X1 U41 ( .A1(n1092), .A2(n380), .ZN(BinLOGIC_25_port) );
  NOR2_X1 U42 ( .A1(n1092), .A2(n377), .ZN(BinLOGIC_30_port) );
  NOR2_X1 U43 ( .A1(n372), .A2(n1092), .ZN(BinLOGIC_12_port) );
  NOR2_X1 U44 ( .A1(n375), .A2(n1092), .ZN(BinLOGIC_10_port) );
  NOR2_X1 U45 ( .A1(n374), .A2(n1091), .ZN(BinLOGIC_11_port) );
  NOR2_X1 U46 ( .A1(n371), .A2(n1091), .ZN(BinLOGIC_5_port) );
  NOR2_X1 U47 ( .A1(n1097), .A2(n371), .ZN(BinMUL_5_port) );
  NOR2_X1 U48 ( .A1(n1098), .A2(n374), .ZN(BinMUL_11_port) );
  OAI22_X1 U49 ( .A1(AorBout_27_port), .A2(n1115), .B1(n570), .B2(n1113), .ZN(
        n92) );
  OAI22_X1 U50 ( .A1(AorBout_26_port), .A2(n1114), .B1(n561), .B2(n1113), .ZN(
        n105) );
  OAI22_X1 U51 ( .A1(AorBout_24_port), .A2(n1115), .B1(n558), .B2(n1113), .ZN(
        n119) );
  OAI22_X1 U52 ( .A1(AorBout_23_port), .A2(n1114), .B1(n562), .B2(n1113), .ZN(
        n126) );
  OAI22_X1 U53 ( .A1(AorBout_22_port), .A2(n1115), .B1(n563), .B2(n1113), .ZN(
        n133) );
  OAI22_X1 U54 ( .A1(AorBout_21_port), .A2(n1114), .B1(n567), .B2(n1113), .ZN(
        n140) );
  OAI22_X1 U55 ( .A1(AorBout_20_port), .A2(n1115), .B1(n559), .B2(n1113), .ZN(
        n147) );
  OAI22_X1 U56 ( .A1(AorBout_30_port), .A2(n1114), .B1(n572), .B2(n1113), .ZN(
        n307) );
  OAI22_X1 U57 ( .A1(AorBout_19_port), .A2(n1115), .B1(n560), .B2(n1112), .ZN(
        n154) );
  OAI22_X1 U58 ( .A1(AorBout_18_port), .A2(n1115), .B1(n564), .B2(n1112), .ZN(
        n161) );
  OAI22_X1 U59 ( .A1(AorBout_17_port), .A2(n1115), .B1(n565), .B2(n1112), .ZN(
        n168) );
  OAI22_X1 U60 ( .A1(AorBout_16_port), .A2(n1115), .B1(n566), .B2(n1112), .ZN(
        n175) );
  OAI22_X1 U61 ( .A1(AorBout_15_port), .A2(n1115), .B1(n549), .B2(n1112), .ZN(
        n182) );
  OAI22_X1 U62 ( .A1(AorBout_14_port), .A2(n1115), .B1(n543), .B2(n1112), .ZN(
        n189) );
  OAI22_X1 U63 ( .A1(AorBout_13_port), .A2(n1115), .B1(n550), .B2(n1112), .ZN(
        n196) );
  OAI22_X1 U64 ( .A1(AorBout_12_port), .A2(n1115), .B1(n544), .B2(n1112), .ZN(
        n203) );
  OAI22_X1 U65 ( .A1(AorBout_11_port), .A2(n1115), .B1(n546), .B2(n1112), .ZN(
        n210) );
  OAI22_X1 U66 ( .A1(AorBout_10_port), .A2(n1115), .B1(n545), .B2(n1112), .ZN(
        n217) );
  OAI22_X1 U67 ( .A1(AorBout_9_port), .A2(n1115), .B1(n551), .B2(n1112), .ZN(
        n224) );
  OAI22_X1 U68 ( .A1(AorBout_8_port), .A2(n1115), .B1(n552), .B2(n1112), .ZN(
        n231) );
  OAI22_X1 U69 ( .A1(AorBout_7_port), .A2(n1114), .B1(n553), .B2(n1112), .ZN(
        n238) );
  OAI22_X1 U70 ( .A1(AorBout_6_port), .A2(n1114), .B1(n554), .B2(n1113), .ZN(
        n245) );
  OAI22_X1 U71 ( .A1(AorBout_5_port), .A2(n1114), .B1(n555), .B2(n1112), .ZN(
        n252) );
  OAI22_X1 U72 ( .A1(AorBout_4_port), .A2(n1114), .B1(n556), .B2(n1113), .ZN(
        n259) );
  OAI22_X1 U73 ( .A1(AorBout_3_port), .A2(n1114), .B1(n557), .B2(n1113), .ZN(
        n266) );
  OAI22_X1 U74 ( .A1(AorBout_2_port), .A2(n1114), .B1(n547), .B2(n1113), .ZN(
        n273) );
  OAI22_X1 U75 ( .A1(AorBout_1_port), .A2(n1114), .B1(n542), .B2(n1113), .ZN(
        n280) );
  OAI22_X1 U76 ( .A1(AorBout_0_port), .A2(n1114), .B1(n548), .B2(n1113), .ZN(
        n287) );
  BUF_X1 U77 ( .A(n87), .Z(n1123) );
  BUF_X1 U78 ( .A(n1069), .Z(n1135) );
  BUF_X1 U79 ( .A(n87), .Z(n1121) );
  BUF_X1 U80 ( .A(n87), .Z(n1122) );
  BUF_X1 U81 ( .A(n98), .Z(n1103) );
  BUF_X1 U82 ( .A(n98), .Z(n1104) );
  NOR2_X1 U83 ( .A1(n1098), .A2(n375), .ZN(BinMUL_10_port) );
  BUF_X1 U84 ( .A(n1069), .Z(n1136) );
  BUF_X1 U85 ( .A(n1069), .Z(n1134) );
  NOR2_X1 U86 ( .A1(n1098), .A2(n372), .ZN(BinMUL_12_port) );
  BUF_X1 U87 ( .A(n98), .Z(n1105) );
  INV_X1 U88 ( .A(n292), .ZN(n1072) );
  INV_X1 U89 ( .A(N1015), .ZN(n96) );
  OR2_X1 U90 ( .A1(n81), .A2(N1020), .ZN(n1076) );
  NOR2_X1 U91 ( .A1(n357), .A2(n1086), .ZN(BinADDSUB_26_port) );
  NOR2_X1 U92 ( .A1(n378), .A2(n1085), .ZN(BinADDSUB_29_port) );
  NOR2_X1 U93 ( .A1(n377), .A2(n1085), .ZN(BinADDSUB_30_port) );
  NOR2_X1 U94 ( .A1(n381), .A2(n1086), .ZN(BinADDSUB_24_port) );
  NOR2_X1 U95 ( .A1(n1088), .A2(n399), .ZN(AinADDSUB_31_port) );
  NOR2_X1 U96 ( .A1(n1087), .A2(n392), .ZN(AinADDSUB_8_port) );
  NOR2_X1 U97 ( .A1(n1087), .A2(n394), .ZN(AinADDSUB_6_port) );
  NOR2_X1 U98 ( .A1(n1087), .A2(n393), .ZN(AinADDSUB_7_port) );
  NOR2_X1 U99 ( .A1(n1089), .A2(n412), .ZN(AinADDSUB_22_port) );
  NOR2_X1 U100 ( .A1(n1088), .A2(n407), .ZN(AinADDSUB_26_port) );
  NOR2_X1 U101 ( .A1(n1088), .A2(n408), .ZN(AinADDSUB_25_port) );
  NOR2_X1 U102 ( .A1(n1088), .A2(n403), .ZN(AinADDSUB_29_port) );
  NOR2_X1 U103 ( .A1(n1089), .A2(n414), .ZN(AinADDSUB_20_port) );
  NOR2_X1 U104 ( .A1(n1088), .A2(n401), .ZN(AinADDSUB_30_port) );
  NOR2_X1 U105 ( .A1(n1089), .A2(n417), .ZN(AinADDSUB_18_port) );
  NOR2_X1 U106 ( .A1(n1088), .A2(n410), .ZN(AinADDSUB_24_port) );
  NOR2_X1 U107 ( .A1(n1089), .A2(n423), .ZN(AinADDSUB_13_port) );
  NOR2_X1 U108 ( .A1(n1089), .A2(n420), .ZN(AinADDSUB_15_port) );
  NOR2_X1 U109 ( .A1(n1089), .A2(n422), .ZN(AinADDSUB_14_port) );
  NOR2_X1 U110 ( .A1(n1089), .A2(n413), .ZN(AinADDSUB_21_port) );
  NOR2_X1 U111 ( .A1(n1089), .A2(n415), .ZN(AinADDSUB_1_port) );
  NOR2_X1 U112 ( .A1(n1089), .A2(n418), .ZN(AinADDSUB_17_port) );
  NOR2_X1 U113 ( .A1(n1088), .A2(n395), .ZN(AinADDSUB_5_port) );
  NOR2_X1 U114 ( .A1(n1089), .A2(n411), .ZN(AinADDSUB_23_port) );
  NOR2_X1 U115 ( .A1(n1089), .A2(n416), .ZN(AinADDSUB_19_port) );
  NOR2_X1 U116 ( .A1(n1088), .A2(n396), .ZN(AinADDSUB_4_port) );
  NOR2_X1 U117 ( .A1(n1089), .A2(n419), .ZN(AinADDSUB_16_port) );
  NOR2_X1 U118 ( .A1(n1090), .A2(n426), .ZN(AinADDSUB_11_port) );
  NOR2_X1 U119 ( .A1(n1090), .A2(n425), .ZN(AinADDSUB_12_port) );
  NOR2_X1 U120 ( .A1(n1090), .A2(n428), .ZN(AinADDSUB_0_port) );
  NOR2_X1 U121 ( .A1(n339), .A2(n1085), .ZN(BinADDSUB_31_port) );
  INV_X1 U122 ( .A(B[5]), .ZN(n371) );
  INV_X1 U123 ( .A(B[24]), .ZN(n381) );
  INV_X1 U124 ( .A(B[30]), .ZN(n377) );
  INV_X1 U125 ( .A(B[29]), .ZN(n378) );
  INV_X1 U126 ( .A(B[23]), .ZN(n383) );
  INV_X1 U127 ( .A(B[18]), .ZN(n384) );
  INV_X1 U128 ( .A(B[25]), .ZN(n380) );
  INV_X1 U129 ( .A(n1078), .ZN(n1116) );
  INV_X1 U130 ( .A(n1077), .ZN(n1114) );
  INV_X1 U131 ( .A(n1079), .ZN(n1112) );
  NOR4_X1 U132 ( .A1(n347), .A2(B[29]), .A3(B[5]), .A4(B[30]), .ZN(n346) );
  NOR2_X1 U133 ( .A1(n1093), .A2(n357), .ZN(BinLOGIC_26_port) );
  NOR2_X1 U134 ( .A1(n1093), .A2(n363), .ZN(BinLOGIC_22_port) );
  NOR2_X1 U135 ( .A1(n1093), .A2(n360), .ZN(BinLOGIC_20_port) );
  NOR2_X1 U136 ( .A1(n1092), .A2(n339), .ZN(BinLOGIC_31_port) );
  NOR2_X1 U137 ( .A1(n1092), .A2(n356), .ZN(BinLOGIC_28_port) );
  NOR2_X1 U138 ( .A1(n1092), .A2(n354), .ZN(BinLOGIC_27_port) );
  NOR2_X1 U139 ( .A1(n1092), .A2(n362), .ZN(BinLOGIC_21_port) );
  BUF_X1 U140 ( .A(n387), .Z(n1088) );
  BUF_X1 U141 ( .A(n387), .Z(n1089) );
  BUF_X1 U142 ( .A(n376), .Z(n1094) );
  BUF_X1 U143 ( .A(n376), .Z(n1095) );
  NOR2_X1 U144 ( .A1(n351), .A2(n1091), .ZN(BinLOGIC_9_port) );
  NOR2_X1 U145 ( .A1(n349), .A2(n1091), .ZN(BinLOGIC_7_port) );
  NOR2_X1 U146 ( .A1(n348), .A2(n1091), .ZN(BinLOGIC_6_port) );
  NOR2_X1 U147 ( .A1(n332), .A2(n1091), .ZN(BinLOGIC_4_port) );
  BUF_X1 U148 ( .A(n376), .Z(n1093) );
  BUF_X1 U149 ( .A(n376), .Z(n1092) );
  NOR2_X1 U150 ( .A1(n1099), .A2(n426), .ZN(AinMUL_11_port) );
  NOR2_X1 U151 ( .A1(n1099), .A2(n398), .ZN(AinMUL_3_port) );
  NOR2_X1 U152 ( .A1(n1098), .A2(n392), .ZN(AinMUL_8_port) );
  NOR2_X1 U153 ( .A1(n1098), .A2(n395), .ZN(AinMUL_5_port) );
  NOR2_X1 U154 ( .A1(n1098), .A2(n428), .ZN(AinMUL_0_port) );
  BUF_X1 U155 ( .A(n376), .Z(n1091) );
  NOR2_X1 U156 ( .A1(n1099), .A2(n420), .ZN(AinMUL_15_port) );
  BUF_X1 U157 ( .A(n90), .Z(n1118) );
  BUF_X1 U158 ( .A(n90), .Z(n1119) );
  BUF_X1 U159 ( .A(n95), .Z(n1109) );
  BUF_X1 U160 ( .A(n95), .Z(n1110) );
  INV_X1 U161 ( .A(n1078), .ZN(n1117) );
  NOR2_X1 U162 ( .A1(n1099), .A2(n415), .ZN(AinMUL_1_port) );
  BUF_X1 U163 ( .A(n99), .Z(n1100) );
  BUF_X1 U164 ( .A(n99), .Z(n1101) );
  INV_X1 U165 ( .A(n1077), .ZN(n1115) );
  NOR2_X1 U166 ( .A1(n1097), .A2(n427), .ZN(AinMUL_10_port) );
  BUF_X1 U167 ( .A(n389), .Z(n1082) );
  BUF_X1 U168 ( .A(n389), .Z(n1083) );
  BUF_X1 U169 ( .A(n369), .Z(n1098) );
  BUF_X1 U170 ( .A(n387), .Z(n1085) );
  BUF_X1 U171 ( .A(n369), .Z(n1099) );
  BUF_X1 U172 ( .A(n389), .Z(n1084) );
  NAND4_X1 U173 ( .A1(n1102), .A2(n1105), .A3(n1078), .A4(n324), .ZN(N1015) );
  NOR4_X1 U174 ( .A1(n1109), .A2(n1118), .A3(n1077), .A4(n1079), .ZN(n324) );
  NOR2_X1 U175 ( .A1(n1094), .A2(n399), .ZN(AinLOGIC_31_port) );
  NOR2_X1 U176 ( .A1(n1094), .A2(n401), .ZN(AinLOGIC_30_port) );
  NOR2_X1 U177 ( .A1(n1094), .A2(n403), .ZN(AinLOGIC_29_port) );
  NOR2_X1 U178 ( .A1(n1094), .A2(n404), .ZN(AinLOGIC_28_port) );
  NOR2_X1 U179 ( .A1(n1094), .A2(n405), .ZN(AinLOGIC_27_port) );
  NOR2_X1 U180 ( .A1(n1094), .A2(n407), .ZN(AinLOGIC_26_port) );
  NOR2_X1 U181 ( .A1(n1094), .A2(n408), .ZN(AinLOGIC_25_port) );
  NOR2_X1 U182 ( .A1(n1095), .A2(n410), .ZN(AinLOGIC_24_port) );
  NOR2_X1 U183 ( .A1(n1095), .A2(n411), .ZN(AinLOGIC_23_port) );
  NOR2_X1 U184 ( .A1(n1095), .A2(n412), .ZN(AinLOGIC_22_port) );
  NOR2_X1 U185 ( .A1(n1095), .A2(n413), .ZN(AinLOGIC_21_port) );
  NOR2_X1 U186 ( .A1(n1095), .A2(n414), .ZN(AinLOGIC_20_port) );
  NOR2_X1 U187 ( .A1(n1095), .A2(n416), .ZN(AinLOGIC_19_port) );
  NOR2_X1 U188 ( .A1(n1095), .A2(n417), .ZN(AinLOGIC_18_port) );
  NOR2_X1 U189 ( .A1(n1095), .A2(n418), .ZN(AinLOGIC_17_port) );
  NOR2_X1 U190 ( .A1(n1095), .A2(n419), .ZN(AinLOGIC_16_port) );
  NOR2_X1 U191 ( .A1(n1095), .A2(n420), .ZN(AinLOGIC_15_port) );
  NOR2_X1 U192 ( .A1(n1095), .A2(n422), .ZN(AinLOGIC_14_port) );
  NOR2_X1 U193 ( .A1(n1094), .A2(n394), .ZN(AinLOGIC_6_port) );
  NOR2_X1 U194 ( .A1(n1094), .A2(n395), .ZN(AinLOGIC_5_port) );
  NOR2_X1 U195 ( .A1(n1094), .A2(n396), .ZN(AinLOGIC_4_port) );
  NOR2_X1 U196 ( .A1(n1094), .A2(n398), .ZN(AinLOGIC_3_port) );
  NOR2_X1 U197 ( .A1(n1094), .A2(n402), .ZN(AinLOGIC_2_port) );
  NOR2_X1 U198 ( .A1(n1095), .A2(n415), .ZN(AinLOGIC_1_port) );
  NOR2_X1 U199 ( .A1(n1096), .A2(n423), .ZN(AinLOGIC_13_port) );
  NOR2_X1 U200 ( .A1(n1096), .A2(n425), .ZN(AinLOGIC_12_port) );
  NOR2_X1 U201 ( .A1(n1096), .A2(n426), .ZN(AinLOGIC_11_port) );
  NOR2_X1 U202 ( .A1(n1096), .A2(n427), .ZN(AinLOGIC_10_port) );
  NOR2_X1 U203 ( .A1(n1093), .A2(n390), .ZN(AinLOGIC_9_port) );
  NOR2_X1 U204 ( .A1(n1093), .A2(n392), .ZN(AinLOGIC_8_port) );
  NOR2_X1 U205 ( .A1(n1093), .A2(n393), .ZN(AinLOGIC_7_port) );
  NOR2_X1 U206 ( .A1(n1092), .A2(n428), .ZN(AinLOGIC_0_port) );
  BUF_X1 U207 ( .A(n387), .Z(n1086) );
  NOR2_X1 U208 ( .A1(n1099), .A2(n422), .ZN(AinMUL_14_port) );
  NOR2_X1 U209 ( .A1(n1099), .A2(n425), .ZN(AinMUL_12_port) );
  NOR2_X1 U210 ( .A1(n1099), .A2(n402), .ZN(AinMUL_2_port) );
  NOR2_X1 U211 ( .A1(n1099), .A2(n423), .ZN(AinMUL_13_port) );
  NOR2_X1 U212 ( .A1(n1097), .A2(n349), .ZN(BinMUL_7_port) );
  NOR2_X1 U213 ( .A1(n332), .A2(n1097), .ZN(BinMUL_4_port) );
  NOR2_X1 U214 ( .A1(n1097), .A2(n348), .ZN(BinMUL_6_port) );
  BUF_X1 U215 ( .A(n95), .Z(n1111) );
  NOR2_X1 U216 ( .A1(n1098), .A2(n393), .ZN(AinMUL_7_port) );
  NOR2_X1 U217 ( .A1(n1098), .A2(n394), .ZN(AinMUL_6_port) );
  NOR2_X1 U218 ( .A1(n1098), .A2(n396), .ZN(AinMUL_4_port) );
  NOR2_X1 U219 ( .A1(n1098), .A2(n390), .ZN(AinMUL_9_port) );
  BUF_X1 U220 ( .A(n369), .Z(n1097) );
  BUF_X1 U221 ( .A(n90), .Z(n1120) );
  BUF_X1 U222 ( .A(n99), .Z(n1102) );
  NOR2_X1 U223 ( .A1(n294), .A2(n289), .ZN(N1021) );
  NOR2_X1 U224 ( .A1(n351), .A2(n1097), .ZN(BinMUL_9_port) );
  AND3_X1 U225 ( .A1(n291), .A2(n329), .A3(n327), .ZN(n1069) );
  NAND4_X1 U226 ( .A1(n292), .A2(n289), .A3(n293), .A4(n294), .ZN(N1008) );
  NOR2_X1 U227 ( .A1(N1019), .A2(N1015), .ZN(n293) );
  AND2_X1 U228 ( .A1(n1111), .A2(n329), .ZN(n87) );
  INV_X1 U229 ( .A(n290), .ZN(N1019) );
  NOR2_X1 U230 ( .A1(n291), .A2(n292), .ZN(N1009) );
  NOR2_X1 U231 ( .A1(n1084), .A2(n398), .ZN(AinSHIFTER_3_port) );
  NOR2_X1 U232 ( .A1(n1084), .A2(n396), .ZN(AinSHIFTER_4_port) );
  NOR2_X1 U233 ( .A1(n1084), .A2(n395), .ZN(AinSHIFTER_5_port) );
  NOR2_X1 U234 ( .A1(n1084), .A2(n394), .ZN(AinSHIFTER_6_port) );
  NOR2_X1 U235 ( .A1(n1084), .A2(n393), .ZN(AinSHIFTER_7_port) );
  NOR2_X1 U236 ( .A1(n1084), .A2(n392), .ZN(AinSHIFTER_8_port) );
  NOR2_X1 U237 ( .A1(n1084), .A2(n390), .ZN(AinSHIFTER_9_port) );
  NOR2_X1 U238 ( .A1(n1084), .A2(n399), .ZN(AinSHIFTER_31_port) );
  INV_X1 U239 ( .A(n294), .ZN(n81) );
  NOR2_X1 U240 ( .A1(n331), .A2(n332), .ZN(Binshift_4_port) );
  NAND2_X1 U241 ( .A1(n295), .A2(n296), .ZN(N1007) );
  AOI22_X1 U242 ( .A1(n1126), .A2(n297), .B1(notAout_31_port), .B2(n1123), 
        .ZN(n296) );
  NAND2_X1 U243 ( .A1(n298), .A2(n299), .ZN(n297) );
  NAND2_X1 U244 ( .A1(n309), .A2(n310), .ZN(N1003) );
  AOI22_X1 U245 ( .A1(n1126), .A2(n311), .B1(notAout_29_port), .B2(n1123), 
        .ZN(n310) );
  NAND2_X1 U246 ( .A1(n312), .A2(n313), .ZN(n311) );
  NAND2_X1 U247 ( .A1(n316), .A2(n317), .ZN(N1001) );
  AOI22_X1 U248 ( .A1(n1124), .A2(n318), .B1(notAout_28_port), .B2(n1123), 
        .ZN(n317) );
  NAND2_X1 U249 ( .A1(n319), .A2(n320), .ZN(n318) );
  NAND2_X1 U250 ( .A1(n107), .A2(n108), .ZN(N995) );
  AOI22_X1 U251 ( .A1(n1124), .A2(n109), .B1(notAout_25_port), .B2(n1121), 
        .ZN(n108) );
  NAND2_X1 U252 ( .A1(n110), .A2(n111), .ZN(n109) );
  NOR2_X1 U253 ( .A1(n1082), .A2(n428), .ZN(AinSHIFTER_0_port) );
  NOR2_X1 U254 ( .A1(n1082), .A2(n415), .ZN(AinSHIFTER_1_port) );
  NOR2_X1 U255 ( .A1(n1083), .A2(n402), .ZN(AinSHIFTER_2_port) );
  NOR2_X1 U256 ( .A1(n1082), .A2(n427), .ZN(AinSHIFTER_10_port) );
  NOR2_X1 U257 ( .A1(n1082), .A2(n426), .ZN(AinSHIFTER_11_port) );
  NOR2_X1 U258 ( .A1(n1082), .A2(n425), .ZN(AinSHIFTER_12_port) );
  NOR2_X1 U259 ( .A1(n1082), .A2(n423), .ZN(AinSHIFTER_13_port) );
  NOR2_X1 U260 ( .A1(n1082), .A2(n422), .ZN(AinSHIFTER_14_port) );
  NOR2_X1 U261 ( .A1(n1082), .A2(n420), .ZN(AinSHIFTER_15_port) );
  NOR2_X1 U262 ( .A1(n1082), .A2(n419), .ZN(AinSHIFTER_16_port) );
  NOR2_X1 U263 ( .A1(n1082), .A2(n418), .ZN(AinSHIFTER_17_port) );
  NOR2_X1 U264 ( .A1(n1082), .A2(n417), .ZN(AinSHIFTER_18_port) );
  NOR2_X1 U265 ( .A1(n1082), .A2(n416), .ZN(AinSHIFTER_19_port) );
  NOR2_X1 U266 ( .A1(n1083), .A2(n414), .ZN(AinSHIFTER_20_port) );
  NOR2_X1 U267 ( .A1(n1083), .A2(n413), .ZN(AinSHIFTER_21_port) );
  NOR2_X1 U268 ( .A1(n1083), .A2(n412), .ZN(AinSHIFTER_22_port) );
  NOR2_X1 U269 ( .A1(n1083), .A2(n411), .ZN(AinSHIFTER_23_port) );
  NOR2_X1 U270 ( .A1(n1083), .A2(n410), .ZN(AinSHIFTER_24_port) );
  NOR2_X1 U271 ( .A1(n1083), .A2(n408), .ZN(AinSHIFTER_25_port) );
  NOR2_X1 U272 ( .A1(n1083), .A2(n407), .ZN(AinSHIFTER_26_port) );
  NOR2_X1 U273 ( .A1(n1083), .A2(n405), .ZN(AinSHIFTER_27_port) );
  NOR2_X1 U274 ( .A1(n1083), .A2(n404), .ZN(AinSHIFTER_28_port) );
  NOR2_X1 U275 ( .A1(n1083), .A2(n403), .ZN(AinSHIFTER_29_port) );
  NOR2_X1 U276 ( .A1(n1083), .A2(n401), .ZN(AinSHIFTER_30_port) );
  NAND2_X1 U277 ( .A1(n83), .A2(n84), .ZN(N999) );
  AOI22_X1 U278 ( .A1(MULout_27_port), .A2(n1134), .B1(ADDSUBout_27_port), 
        .B2(n1131), .ZN(n83) );
  AOI22_X1 U279 ( .A1(n1125), .A2(n86), .B1(notAout_27_port), .B2(n1121), .ZN(
        n84) );
  NAND2_X1 U280 ( .A1(n100), .A2(n101), .ZN(N997) );
  AOI22_X1 U281 ( .A1(MULout_26_port), .A2(n1134), .B1(ADDSUBout_26_port), 
        .B2(n1131), .ZN(n100) );
  AOI22_X1 U282 ( .A1(n1124), .A2(n102), .B1(notAout_26_port), .B2(n1121), 
        .ZN(n101) );
  NAND2_X1 U283 ( .A1(n114), .A2(n115), .ZN(N993) );
  AOI22_X1 U284 ( .A1(MULout_24_port), .A2(n1134), .B1(ADDSUBout_24_port), 
        .B2(n1131), .ZN(n114) );
  AOI22_X1 U285 ( .A1(n1124), .A2(n116), .B1(notAout_24_port), .B2(n1121), 
        .ZN(n115) );
  NAND2_X1 U286 ( .A1(n121), .A2(n122), .ZN(N991) );
  AOI22_X1 U287 ( .A1(MULout_23_port), .A2(n1134), .B1(ADDSUBout_23_port), 
        .B2(n1131), .ZN(n121) );
  AOI22_X1 U288 ( .A1(n1124), .A2(n123), .B1(notAout_23_port), .B2(n1121), 
        .ZN(n122) );
  NAND2_X1 U289 ( .A1(n128), .A2(n129), .ZN(N989) );
  AOI22_X1 U290 ( .A1(MULout_22_port), .A2(n1134), .B1(ADDSUBout_22_port), 
        .B2(n1131), .ZN(n128) );
  AOI22_X1 U291 ( .A1(n1124), .A2(n130), .B1(notAout_22_port), .B2(n1121), 
        .ZN(n129) );
  NAND2_X1 U292 ( .A1(n135), .A2(n136), .ZN(N987) );
  AOI22_X1 U293 ( .A1(MULout_21_port), .A2(n1134), .B1(ADDSUBout_21_port), 
        .B2(n1131), .ZN(n135) );
  AOI22_X1 U294 ( .A1(n1124), .A2(n137), .B1(notAout_21_port), .B2(n1121), 
        .ZN(n136) );
  NAND2_X1 U295 ( .A1(n142), .A2(n143), .ZN(N985) );
  AOI22_X1 U296 ( .A1(MULout_20_port), .A2(n1135), .B1(ADDSUBout_20_port), 
        .B2(n1132), .ZN(n142) );
  AOI22_X1 U297 ( .A1(n1124), .A2(n144), .B1(notAout_20_port), .B2(n1121), 
        .ZN(n143) );
  NAND2_X1 U298 ( .A1(n149), .A2(n150), .ZN(N983) );
  AOI22_X1 U299 ( .A1(MULout_19_port), .A2(n1134), .B1(ADDSUBout_19_port), 
        .B2(n1131), .ZN(n149) );
  AOI22_X1 U300 ( .A1(n1124), .A2(n151), .B1(notAout_19_port), .B2(n1121), 
        .ZN(n150) );
  NAND2_X1 U301 ( .A1(n156), .A2(n157), .ZN(N981) );
  AOI22_X1 U302 ( .A1(MULout_18_port), .A2(n1134), .B1(ADDSUBout_18_port), 
        .B2(n1131), .ZN(n156) );
  AOI22_X1 U303 ( .A1(n1124), .A2(n158), .B1(notAout_18_port), .B2(n1121), 
        .ZN(n157) );
  NAND2_X1 U304 ( .A1(n163), .A2(n164), .ZN(N979) );
  AOI22_X1 U305 ( .A1(MULout_17_port), .A2(n1134), .B1(ADDSUBout_17_port), 
        .B2(n1131), .ZN(n163) );
  AOI22_X1 U306 ( .A1(n1124), .A2(n165), .B1(notAout_17_port), .B2(n1121), 
        .ZN(n164) );
  NAND2_X1 U307 ( .A1(n170), .A2(n171), .ZN(N977) );
  AOI22_X1 U308 ( .A1(MULout_16_port), .A2(n1134), .B1(ADDSUBout_16_port), 
        .B2(n1132), .ZN(n170) );
  AOI22_X1 U309 ( .A1(n1124), .A2(n172), .B1(notAout_16_port), .B2(n1121), 
        .ZN(n171) );
  NAND2_X1 U310 ( .A1(n177), .A2(n178), .ZN(N975) );
  AOI22_X1 U311 ( .A1(MULout_15_port), .A2(n1135), .B1(ADDSUBout_15_port), 
        .B2(n1132), .ZN(n177) );
  AOI22_X1 U312 ( .A1(n1125), .A2(n179), .B1(notAout_15_port), .B2(n1122), 
        .ZN(n178) );
  NAND2_X1 U313 ( .A1(n184), .A2(n185), .ZN(N973) );
  AOI22_X1 U314 ( .A1(MULout_14_port), .A2(n1135), .B1(ADDSUBout_14_port), 
        .B2(n1132), .ZN(n184) );
  AOI22_X1 U315 ( .A1(n1125), .A2(n186), .B1(notAout_14_port), .B2(n1122), 
        .ZN(n185) );
  NAND2_X1 U316 ( .A1(n191), .A2(n192), .ZN(N971) );
  AOI22_X1 U317 ( .A1(MULout_13_port), .A2(n1135), .B1(ADDSUBout_13_port), 
        .B2(n1132), .ZN(n191) );
  AOI22_X1 U318 ( .A1(n1125), .A2(n193), .B1(notAout_13_port), .B2(n1122), 
        .ZN(n192) );
  NAND2_X1 U319 ( .A1(n198), .A2(n199), .ZN(N969) );
  AOI22_X1 U320 ( .A1(MULout_12_port), .A2(n1135), .B1(ADDSUBout_12_port), 
        .B2(n1132), .ZN(n198) );
  AOI22_X1 U321 ( .A1(n1125), .A2(n200), .B1(notAout_12_port), .B2(n1122), 
        .ZN(n199) );
  NAND2_X1 U322 ( .A1(n205), .A2(n206), .ZN(N967) );
  AOI22_X1 U323 ( .A1(MULout_11_port), .A2(n1135), .B1(ADDSUBout_11_port), 
        .B2(n1132), .ZN(n205) );
  AOI22_X1 U324 ( .A1(n1125), .A2(n207), .B1(notAout_11_port), .B2(n1122), 
        .ZN(n206) );
  NAND2_X1 U325 ( .A1(n212), .A2(n213), .ZN(N965) );
  AOI22_X1 U326 ( .A1(MULout_10_port), .A2(n1135), .B1(ADDSUBout_10_port), 
        .B2(n1132), .ZN(n212) );
  AOI22_X1 U327 ( .A1(n1125), .A2(n214), .B1(notAout_10_port), .B2(n1122), 
        .ZN(n213) );
  NAND2_X1 U328 ( .A1(n219), .A2(n220), .ZN(N963) );
  AOI22_X1 U329 ( .A1(MULout_9_port), .A2(n1135), .B1(ADDSUBout_9_port), .B2(
        n1132), .ZN(n219) );
  AOI22_X1 U330 ( .A1(n1125), .A2(n221), .B1(notAout_9_port), .B2(n1122), .ZN(
        n220) );
  NAND2_X1 U331 ( .A1(n226), .A2(n227), .ZN(N961) );
  AOI22_X1 U332 ( .A1(MULout_8_port), .A2(n1135), .B1(ADDSUBout_8_port), .B2(
        n1132), .ZN(n226) );
  AOI22_X1 U333 ( .A1(n1125), .A2(n228), .B1(notAout_8_port), .B2(n1122), .ZN(
        n227) );
  NAND2_X1 U334 ( .A1(n233), .A2(n234), .ZN(N959) );
  AOI22_X1 U335 ( .A1(MULout_7_port), .A2(n1135), .B1(ADDSUBout_7_port), .B2(
        n1132), .ZN(n233) );
  AOI22_X1 U336 ( .A1(n1125), .A2(n235), .B1(notAout_7_port), .B2(n1122), .ZN(
        n234) );
  NAND2_X1 U337 ( .A1(n240), .A2(n241), .ZN(N957) );
  AOI22_X1 U338 ( .A1(MULout_6_port), .A2(n1135), .B1(ADDSUBout_6_port), .B2(
        n1132), .ZN(n240) );
  AOI22_X1 U339 ( .A1(n1125), .A2(n242), .B1(notAout_6_port), .B2(n1122), .ZN(
        n241) );
  NAND2_X1 U340 ( .A1(n247), .A2(n248), .ZN(N955) );
  AOI22_X1 U341 ( .A1(MULout_5_port), .A2(n1135), .B1(ADDSUBout_5_port), .B2(
        n1133), .ZN(n247) );
  AOI22_X1 U342 ( .A1(n1125), .A2(n249), .B1(notAout_5_port), .B2(n1122), .ZN(
        n248) );
  NAND2_X1 U343 ( .A1(n302), .A2(n303), .ZN(N1005) );
  AOI22_X1 U344 ( .A1(MULout_30_port), .A2(n1136), .B1(ADDSUBout_30_port), 
        .B2(n1133), .ZN(n302) );
  AOI22_X1 U345 ( .A1(n1126), .A2(n304), .B1(notAout_30_port), .B2(n1123), 
        .ZN(n303) );
  NAND2_X1 U346 ( .A1(n254), .A2(n255), .ZN(N953) );
  AOI22_X1 U347 ( .A1(MULout_4_port), .A2(n1136), .B1(ADDSUBout_4_port), .B2(
        n1133), .ZN(n254) );
  AOI22_X1 U348 ( .A1(n1126), .A2(n256), .B1(notAout_4_port), .B2(n1122), .ZN(
        n255) );
  NAND2_X1 U349 ( .A1(n261), .A2(n262), .ZN(N951) );
  AOI22_X1 U350 ( .A1(MULout_3_port), .A2(n1136), .B1(ADDSUBout_3_port), .B2(
        n1133), .ZN(n261) );
  AOI22_X1 U351 ( .A1(n1126), .A2(n263), .B1(notAout_3_port), .B2(n1123), .ZN(
        n262) );
  NAND2_X1 U352 ( .A1(n268), .A2(n269), .ZN(N949) );
  AOI22_X1 U353 ( .A1(MULout_2_port), .A2(n1136), .B1(ADDSUBout_2_port), .B2(
        n1133), .ZN(n268) );
  AOI22_X1 U354 ( .A1(n1126), .A2(n270), .B1(notAout_2_port), .B2(n1123), .ZN(
        n269) );
  NAND2_X1 U355 ( .A1(n275), .A2(n276), .ZN(N947) );
  AOI22_X1 U356 ( .A1(MULout_1_port), .A2(n1136), .B1(ADDSUBout_1_port), .B2(
        n1133), .ZN(n275) );
  AOI22_X1 U357 ( .A1(n1126), .A2(n277), .B1(notAout_1_port), .B2(n1123), .ZN(
        n276) );
  NAND2_X1 U358 ( .A1(n282), .A2(n283), .ZN(N945) );
  AOI22_X1 U359 ( .A1(MULout_0_port), .A2(n1136), .B1(ADDSUBout_0_port), .B2(
        n1133), .ZN(n282) );
  AOI22_X1 U360 ( .A1(n1126), .A2(n284), .B1(notAout_0_port), .B2(n1123), .ZN(
        n283) );
  INV_X1 U361 ( .A(n82), .ZN(complete) );
  INV_X1 U362 ( .A(A[0]), .ZN(n428) );
  INV_X1 U363 ( .A(A[12]), .ZN(n425) );
  INV_X1 U364 ( .A(A[8]), .ZN(n392) );
  INV_X1 U365 ( .A(A[1]), .ZN(n415) );
  INV_X1 U366 ( .A(A[7]), .ZN(n393) );
  INV_X1 U367 ( .A(A[5]), .ZN(n395) );
  INV_X1 U368 ( .A(A[6]), .ZN(n394) );
  INV_X1 U369 ( .A(A[4]), .ZN(n396) );
  INV_X1 U370 ( .A(B[4]), .ZN(n332) );
  INV_X1 U371 ( .A(B[9]), .ZN(n351) );
  INV_X1 U372 ( .A(B[7]), .ZN(n349) );
  INV_X1 U373 ( .A(B[6]), .ZN(n348) );
  INV_X1 U374 ( .A(A[31]), .ZN(n399) );
  INV_X1 U375 ( .A(A[26]), .ZN(n407) );
  INV_X1 U376 ( .A(A[25]), .ZN(n408) );
  INV_X1 U377 ( .A(A[27]), .ZN(n405) );
  INV_X1 U378 ( .A(A[28]), .ZN(n404) );
  INV_X1 U379 ( .A(A[24]), .ZN(n410) );
  INV_X1 U380 ( .A(A[20]), .ZN(n414) );
  INV_X1 U381 ( .A(A[22]), .ZN(n412) );
  INV_X1 U382 ( .A(A[18]), .ZN(n417) );
  INV_X1 U383 ( .A(A[21]), .ZN(n413) );
  INV_X1 U384 ( .A(A[17]), .ZN(n418) );
  INV_X1 U385 ( .A(A[23]), .ZN(n411) );
  INV_X1 U386 ( .A(A[19]), .ZN(n416) );
  INV_X1 U387 ( .A(A[16]), .ZN(n419) );
  INV_X1 U388 ( .A(B[26]), .ZN(n357) );
  INV_X1 U389 ( .A(B[14]), .ZN(n366) );
  INV_X1 U390 ( .A(B[8]), .ZN(n350) );
  INV_X1 U391 ( .A(B[21]), .ZN(n362) );
  INV_X1 U392 ( .A(B[20]), .ZN(n360) );
  INV_X1 U393 ( .A(B[31]), .ZN(n339) );
  INV_X1 U394 ( .A(A[29]), .ZN(n403) );
  INV_X1 U395 ( .A(A[30]), .ZN(n401) );
  NOR3_X1 U396 ( .A1(ALUsel[0]), .A2(ALUsel[3]), .A3(n289), .ZN(n90) );
  AOI221_X1 U397 ( .B1(AxorBout_31_port), .B2(n1111), .C1(SHIFTERout_31_port), 
        .C2(n1108), .A(n301), .ZN(n298) );
  OAI22_X1 U398 ( .A1(n345), .A2(n1105), .B1(AxorBout_31_port), .B2(n1102), 
        .ZN(n301) );
  AOI221_X1 U399 ( .B1(AxorBout_29_port), .B2(n1111), .C1(SHIFTERout_29_port), 
        .C2(n1108), .A(n315), .ZN(n312) );
  OAI22_X1 U400 ( .A1(n391), .A2(n1105), .B1(AxorBout_29_port), .B2(n1102), 
        .ZN(n315) );
  AOI221_X1 U401 ( .B1(AxorBout_28_port), .B2(n1111), .C1(SHIFTERout_28_port), 
        .C2(n1106), .A(n322), .ZN(n319) );
  OAI22_X1 U402 ( .A1(n352), .A2(n1105), .B1(AxorBout_28_port), .B2(n1102), 
        .ZN(n322) );
  AOI221_X1 U403 ( .B1(AxorBout_25_port), .B2(n1109), .C1(SHIFTERout_25_port), 
        .C2(n1106), .A(n113), .ZN(n110) );
  OAI22_X1 U404 ( .A1(n373), .A2(n1103), .B1(AxorBout_25_port), .B2(n1100), 
        .ZN(n113) );
  NAND2_X1 U405 ( .A1(ALUsel[2]), .A2(n328), .ZN(n289) );
  INV_X1 U406 ( .A(ALUsel[1]), .ZN(n328) );
  INV_X1 U407 ( .A(ALUsel[0]), .ZN(n291) );
  NAND4_X1 U408 ( .A1(enSHIFTER), .A2(n338), .A3(N1019), .A4(n339), .ZN(n82)
         );
  NAND4_X1 U409 ( .A1(n341), .A2(n343), .A3(n344), .A4(n346), .ZN(n338) );
  NOR4_X1 U410 ( .A1(n358), .A2(B[16]), .A3(B[18]), .A4(B[17]), .ZN(n343) );
  NOR4_X1 U411 ( .A1(n353), .A2(B[23]), .A3(B[25]), .A4(B[24]), .ZN(n344) );
  NOR2_X1 U412 ( .A1(n328), .A2(ALUsel[3]), .ZN(n327) );
  AND4_X1 U413 ( .A1(ALUsel[0]), .A2(ALUsel[3]), .A3(n328), .A4(n329), .ZN(
        n1077) );
  OR3_X1 U414 ( .A1(n291), .A2(ALUsel[3]), .A3(n289), .ZN(n1078) );
  NAND2_X1 U415 ( .A1(enSHIFTER), .A2(n82), .ZN(n331) );
  NOR2_X1 U416 ( .A1(n340), .A2(N1021), .ZN(n290) );
  NOR4_X1 U417 ( .A1(n291), .A2(n328), .A3(n330), .A4(ALUsel[2]), .ZN(n340) );
  INV_X1 U418 ( .A(ALUsel[2]), .ZN(n329) );
  NAND2_X1 U419 ( .A1(ALUsel[3]), .A2(n291), .ZN(n294) );
  AND3_X1 U420 ( .A1(n327), .A2(n291), .A3(ALUsel[2]), .ZN(n1079) );
  INV_X1 U421 ( .A(enADDSUB), .ZN(n387) );
  INV_X1 U422 ( .A(enLOGIC), .ZN(n376) );
  AND2_X1 U423 ( .A1(ALUsel[0]), .A2(n327), .ZN(n95) );
  INV_X1 U424 ( .A(enSHIFTER), .ZN(n389) );
  NAND2_X1 U425 ( .A1(n305), .A2(n306), .ZN(n304) );
  AOI221_X1 U426 ( .B1(AxorBout_30_port), .B2(n1111), .C1(SHIFTERout_30_port), 
        .C2(n1108), .A(n308), .ZN(n305) );
  AOI221_X1 U427 ( .B1(notBout_30_port), .B2(n1118), .C1(n388), .C2(n1116), 
        .A(n307), .ZN(n306) );
  OAI22_X1 U428 ( .A1(n388), .A2(n1105), .B1(AxorBout_30_port), .B2(n1102), 
        .ZN(n308) );
  NAND2_X1 U429 ( .A1(n271), .A2(n272), .ZN(n270) );
  AOI221_X1 U430 ( .B1(AxorBout_2_port), .B2(n1111), .C1(SHIFTERout_2_port), 
        .C2(n1108), .A(n274), .ZN(n271) );
  AOI221_X1 U431 ( .B1(notBout_2_port), .B2(n1118), .C1(n397), .C2(n1116), .A(
        n273), .ZN(n272) );
  OAI22_X1 U432 ( .A1(n397), .A2(n1105), .B1(AxorBout_2_port), .B2(n1102), 
        .ZN(n274) );
  NAND2_X1 U433 ( .A1(n278), .A2(n279), .ZN(n277) );
  AOI221_X1 U434 ( .B1(AxorBout_1_port), .B2(n1111), .C1(SHIFTERout_1_port), 
        .C2(n1108), .A(n281), .ZN(n278) );
  AOI221_X1 U435 ( .B1(notBout_1_port), .B2(n1118), .C1(n400), .C2(n1116), .A(
        n280), .ZN(n279) );
  OAI22_X1 U436 ( .A1(n400), .A2(n1105), .B1(AxorBout_1_port), .B2(n1102), 
        .ZN(n281) );
  NAND2_X1 U437 ( .A1(n285), .A2(n286), .ZN(n284) );
  AOI221_X1 U438 ( .B1(AxorBout_0_port), .B2(n1111), .C1(SHIFTERout_0_port), 
        .C2(n1108), .A(n288), .ZN(n285) );
  AOI221_X1 U439 ( .B1(notBout_0_port), .B2(n1118), .C1(n455), .C2(n1116), .A(
        n287), .ZN(n286) );
  OAI22_X1 U440 ( .A1(n455), .A2(n1105), .B1(AxorBout_0_port), .B2(n1102), 
        .ZN(n288) );
  NAND2_X1 U441 ( .A1(n88), .A2(n89), .ZN(n86) );
  AOI221_X1 U442 ( .B1(AxorBout_27_port), .B2(n1110), .C1(SHIFTERout_27_port), 
        .C2(n1107), .A(n97), .ZN(n88) );
  AOI221_X1 U443 ( .B1(notBout_27_port), .B2(n1120), .C1(n364), .C2(n1117), 
        .A(n92), .ZN(n89) );
  OAI22_X1 U444 ( .A1(n364), .A2(n1103), .B1(AxorBout_27_port), .B2(n1100), 
        .ZN(n97) );
  NAND2_X1 U445 ( .A1(n103), .A2(n104), .ZN(n102) );
  AOI221_X1 U446 ( .B1(AxorBout_26_port), .B2(n1109), .C1(SHIFTERout_26_port), 
        .C2(n1106), .A(n106), .ZN(n103) );
  AOI221_X1 U447 ( .B1(notBout_26_port), .B2(n1120), .C1(n370), .C2(n1116), 
        .A(n105), .ZN(n104) );
  OAI22_X1 U448 ( .A1(n370), .A2(n1103), .B1(AxorBout_26_port), .B2(n1100), 
        .ZN(n106) );
  NAND2_X1 U449 ( .A1(n117), .A2(n118), .ZN(n116) );
  AOI221_X1 U450 ( .B1(AxorBout_24_port), .B2(n1109), .C1(SHIFTERout_24_port), 
        .C2(n1106), .A(n120), .ZN(n117) );
  AOI221_X1 U451 ( .B1(notBout_24_port), .B2(n1120), .C1(n336), .C2(n1117), 
        .A(n119), .ZN(n118) );
  OAI22_X1 U452 ( .A1(n336), .A2(n1103), .B1(AxorBout_24_port), .B2(n1100), 
        .ZN(n120) );
  NAND2_X1 U453 ( .A1(n124), .A2(n125), .ZN(n123) );
  AOI221_X1 U454 ( .B1(AxorBout_23_port), .B2(n1109), .C1(SHIFTERout_23_port), 
        .C2(n1106), .A(n127), .ZN(n124) );
  AOI221_X1 U455 ( .B1(notBout_23_port), .B2(n1120), .C1(n379), .C2(n1116), 
        .A(n126), .ZN(n125) );
  OAI22_X1 U456 ( .A1(n379), .A2(n1103), .B1(AxorBout_23_port), .B2(n1100), 
        .ZN(n127) );
  NAND2_X1 U457 ( .A1(n131), .A2(n132), .ZN(n130) );
  AOI221_X1 U458 ( .B1(AxorBout_22_port), .B2(n1109), .C1(SHIFTERout_22_port), 
        .C2(n1106), .A(n134), .ZN(n131) );
  AOI221_X1 U459 ( .B1(notBout_22_port), .B2(n1120), .C1(n382), .C2(n1117), 
        .A(n133), .ZN(n132) );
  OAI22_X1 U460 ( .A1(n382), .A2(n1103), .B1(AxorBout_22_port), .B2(n1100), 
        .ZN(n134) );
  NAND2_X1 U461 ( .A1(n138), .A2(n139), .ZN(n137) );
  AOI221_X1 U462 ( .B1(AxorBout_21_port), .B2(n1109), .C1(SHIFTERout_21_port), 
        .C2(n1106), .A(n141), .ZN(n138) );
  AOI221_X1 U463 ( .B1(notBout_21_port), .B2(n1120), .C1(n342), .C2(n1116), 
        .A(n140), .ZN(n139) );
  OAI22_X1 U464 ( .A1(n342), .A2(n1103), .B1(AxorBout_21_port), .B2(n1100), 
        .ZN(n141) );
  NAND2_X1 U465 ( .A1(n145), .A2(n146), .ZN(n144) );
  AOI221_X1 U466 ( .B1(AxorBout_20_port), .B2(n1109), .C1(SHIFTERout_20_port), 
        .C2(n1106), .A(n148), .ZN(n145) );
  AOI221_X1 U467 ( .B1(notBout_20_port), .B2(n1119), .C1(n355), .C2(n1117), 
        .A(n147), .ZN(n146) );
  OAI22_X1 U468 ( .A1(n355), .A2(n1103), .B1(AxorBout_20_port), .B2(n1100), 
        .ZN(n148) );
  NAND2_X1 U469 ( .A1(n152), .A2(n153), .ZN(n151) );
  AOI221_X1 U470 ( .B1(AxorBout_19_port), .B2(n1109), .C1(SHIFTERout_19_port), 
        .C2(n1106), .A(n155), .ZN(n152) );
  AOI221_X1 U471 ( .B1(notBout_19_port), .B2(n1119), .C1(n361), .C2(n1117), 
        .A(n154), .ZN(n153) );
  OAI22_X1 U472 ( .A1(n361), .A2(n1103), .B1(AxorBout_19_port), .B2(n1100), 
        .ZN(n155) );
  NAND2_X1 U473 ( .A1(n159), .A2(n160), .ZN(n158) );
  AOI221_X1 U474 ( .B1(AxorBout_18_port), .B2(n1109), .C1(SHIFTERout_18_port), 
        .C2(n1106), .A(n162), .ZN(n159) );
  AOI221_X1 U475 ( .B1(notBout_18_port), .B2(n1119), .C1(n406), .C2(n1117), 
        .A(n161), .ZN(n160) );
  OAI22_X1 U476 ( .A1(n406), .A2(n1103), .B1(AxorBout_18_port), .B2(n1100), 
        .ZN(n162) );
  NAND2_X1 U477 ( .A1(n166), .A2(n167), .ZN(n165) );
  AOI221_X1 U478 ( .B1(AxorBout_17_port), .B2(n1109), .C1(SHIFTERout_17_port), 
        .C2(n1106), .A(n169), .ZN(n166) );
  AOI221_X1 U479 ( .B1(notBout_17_port), .B2(n1119), .C1(n409), .C2(n1117), 
        .A(n168), .ZN(n167) );
  OAI22_X1 U480 ( .A1(n409), .A2(n1103), .B1(AxorBout_17_port), .B2(n1100), 
        .ZN(n169) );
  NAND2_X1 U481 ( .A1(n173), .A2(n174), .ZN(n172) );
  AOI221_X1 U482 ( .B1(AxorBout_16_port), .B2(n1109), .C1(SHIFTERout_16_port), 
        .C2(n1106), .A(n176), .ZN(n173) );
  AOI221_X1 U483 ( .B1(notBout_16_port), .B2(n1119), .C1(n421), .C2(n1117), 
        .A(n175), .ZN(n174) );
  OAI22_X1 U484 ( .A1(n421), .A2(n1103), .B1(AxorBout_16_port), .B2(n1100), 
        .ZN(n176) );
  NAND2_X1 U485 ( .A1(n180), .A2(n181), .ZN(n179) );
  AOI221_X1 U486 ( .B1(AxorBout_15_port), .B2(n1109), .C1(SHIFTERout_15_port), 
        .C2(n1107), .A(n183), .ZN(n180) );
  AOI221_X1 U487 ( .B1(notBout_15_port), .B2(n1119), .C1(n424), .C2(n1117), 
        .A(n182), .ZN(n181) );
  OAI22_X1 U488 ( .A1(n424), .A2(n1104), .B1(AxorBout_15_port), .B2(n1101), 
        .ZN(n183) );
  NAND2_X1 U489 ( .A1(n187), .A2(n188), .ZN(n186) );
  AOI221_X1 U490 ( .B1(AxorBout_14_port), .B2(n1110), .C1(SHIFTERout_14_port), 
        .C2(n1107), .A(n190), .ZN(n187) );
  AOI221_X1 U491 ( .B1(notBout_14_port), .B2(n1119), .C1(n430), .C2(n1117), 
        .A(n189), .ZN(n188) );
  OAI22_X1 U492 ( .A1(n430), .A2(n1104), .B1(AxorBout_14_port), .B2(n1101), 
        .ZN(n190) );
  NAND2_X1 U493 ( .A1(n194), .A2(n195), .ZN(n193) );
  AOI221_X1 U494 ( .B1(AxorBout_13_port), .B2(n1110), .C1(SHIFTERout_13_port), 
        .C2(n1107), .A(n197), .ZN(n194) );
  AOI221_X1 U495 ( .B1(notBout_13_port), .B2(n1119), .C1(n539), .C2(n1117), 
        .A(n196), .ZN(n195) );
  OAI22_X1 U496 ( .A1(n539), .A2(n1104), .B1(AxorBout_13_port), .B2(n1101), 
        .ZN(n197) );
  NAND2_X1 U497 ( .A1(n201), .A2(n202), .ZN(n200) );
  AOI221_X1 U498 ( .B1(AxorBout_12_port), .B2(n1110), .C1(SHIFTERout_12_port), 
        .C2(n1107), .A(n204), .ZN(n201) );
  AOI221_X1 U499 ( .B1(notBout_12_port), .B2(n1119), .C1(n540), .C2(n1117), 
        .A(n203), .ZN(n202) );
  OAI22_X1 U500 ( .A1(n540), .A2(n1104), .B1(AxorBout_12_port), .B2(n1101), 
        .ZN(n204) );
  NAND2_X1 U501 ( .A1(n208), .A2(n209), .ZN(n207) );
  AOI221_X1 U502 ( .B1(AxorBout_11_port), .B2(n1110), .C1(SHIFTERout_11_port), 
        .C2(n1107), .A(n211), .ZN(n208) );
  AOI221_X1 U503 ( .B1(notBout_11_port), .B2(n1119), .C1(n538), .C2(n1117), 
        .A(n210), .ZN(n209) );
  OAI22_X1 U504 ( .A1(n538), .A2(n1104), .B1(AxorBout_11_port), .B2(n1101), 
        .ZN(n211) );
  NAND2_X1 U505 ( .A1(n215), .A2(n216), .ZN(n214) );
  AOI221_X1 U506 ( .B1(AxorBout_10_port), .B2(n1110), .C1(SHIFTERout_10_port), 
        .C2(n1107), .A(n218), .ZN(n215) );
  AOI221_X1 U507 ( .B1(notBout_10_port), .B2(n1119), .C1(n541), .C2(n1117), 
        .A(n217), .ZN(n216) );
  OAI22_X1 U508 ( .A1(n541), .A2(n1104), .B1(AxorBout_10_port), .B2(n1101), 
        .ZN(n218) );
  NAND2_X1 U509 ( .A1(n222), .A2(n223), .ZN(n221) );
  AOI221_X1 U510 ( .B1(AxorBout_9_port), .B2(n1110), .C1(SHIFTERout_9_port), 
        .C2(n1107), .A(n225), .ZN(n222) );
  AOI221_X1 U511 ( .B1(notBout_9_port), .B2(n1119), .C1(n433), .C2(n1117), .A(
        n224), .ZN(n223) );
  OAI22_X1 U512 ( .A1(n433), .A2(n1104), .B1(AxorBout_9_port), .B2(n1101), 
        .ZN(n225) );
  NAND2_X1 U513 ( .A1(n229), .A2(n230), .ZN(n228) );
  AOI221_X1 U514 ( .B1(AxorBout_8_port), .B2(n1110), .C1(SHIFTERout_8_port), 
        .C2(n1107), .A(n232), .ZN(n229) );
  AOI221_X1 U515 ( .B1(notBout_8_port), .B2(n1119), .C1(n439), .C2(n1117), .A(
        n231), .ZN(n230) );
  OAI22_X1 U516 ( .A1(n439), .A2(n1104), .B1(AxorBout_8_port), .B2(n1101), 
        .ZN(n232) );
  NAND2_X1 U517 ( .A1(n236), .A2(n237), .ZN(n235) );
  AOI221_X1 U518 ( .B1(AxorBout_7_port), .B2(n1110), .C1(SHIFTERout_7_port), 
        .C2(n1107), .A(n239), .ZN(n236) );
  AOI221_X1 U519 ( .B1(notBout_7_port), .B2(n1118), .C1(n442), .C2(n1116), .A(
        n238), .ZN(n237) );
  OAI22_X1 U520 ( .A1(n442), .A2(n1104), .B1(AxorBout_7_port), .B2(n1101), 
        .ZN(n239) );
  NAND2_X1 U521 ( .A1(n243), .A2(n244), .ZN(n242) );
  AOI221_X1 U522 ( .B1(AxorBout_6_port), .B2(n1110), .C1(SHIFTERout_6_port), 
        .C2(n1107), .A(n246), .ZN(n243) );
  AOI221_X1 U523 ( .B1(notBout_6_port), .B2(n1118), .C1(n448), .C2(n1116), .A(
        n245), .ZN(n244) );
  OAI22_X1 U524 ( .A1(n448), .A2(n1104), .B1(AxorBout_6_port), .B2(n1101), 
        .ZN(n246) );
  NAND2_X1 U525 ( .A1(n250), .A2(n251), .ZN(n249) );
  AOI221_X1 U526 ( .B1(AxorBout_5_port), .B2(n1110), .C1(SHIFTERout_5_port), 
        .C2(n1107), .A(n253), .ZN(n250) );
  AOI221_X1 U527 ( .B1(notBout_5_port), .B2(n1118), .C1(n451), .C2(n1116), .A(
        n252), .ZN(n251) );
  OAI22_X1 U528 ( .A1(n451), .A2(n1104), .B1(AxorBout_5_port), .B2(n1101), 
        .ZN(n253) );
  NAND2_X1 U529 ( .A1(n257), .A2(n258), .ZN(n256) );
  AOI221_X1 U530 ( .B1(AxorBout_4_port), .B2(n1110), .C1(SHIFTERout_4_port), 
        .C2(n1108), .A(n260), .ZN(n257) );
  AOI221_X1 U531 ( .B1(notBout_4_port), .B2(n1118), .C1(n452), .C2(n1116), .A(
        n259), .ZN(n258) );
  OAI22_X1 U532 ( .A1(n452), .A2(n1104), .B1(AxorBout_4_port), .B2(n1101), 
        .ZN(n260) );
  NAND2_X1 U533 ( .A1(n264), .A2(n265), .ZN(n263) );
  AOI221_X1 U534 ( .B1(AxorBout_3_port), .B2(n1110), .C1(SHIFTERout_3_port), 
        .C2(n1108), .A(n267), .ZN(n264) );
  AOI221_X1 U535 ( .B1(notBout_3_port), .B2(n1118), .C1(n454), .C2(n1116), .A(
        n266), .ZN(n265) );
  OAI22_X1 U536 ( .A1(n454), .A2(n1105), .B1(AxorBout_3_port), .B2(n1102), 
        .ZN(n267) );
  INV_X1 U537 ( .A(enMUL), .ZN(n369) );
  INV_X1 U538 ( .A(ALUsel[3]), .ZN(n330) );
  NOR2_X1 U539 ( .A1(n380), .A2(n1086), .ZN(BinADDSUB_25_port) );
  NOR2_X1 U540 ( .A1(n384), .A2(n1086), .ZN(BinADDSUB_18_port) );
  NOR2_X1 U541 ( .A1(n363), .A2(n1086), .ZN(BinADDSUB_22_port) );
  INV_X1 U542 ( .A(B[22]), .ZN(n363) );
  INV_X1 U543 ( .A(B[13]), .ZN(n368) );
  NOR2_X1 U544 ( .A1(n333), .A2(n1091), .ZN(BinLOGIC_3_port) );
  NOR2_X1 U545 ( .A1(n333), .A2(n1097), .ZN(BinMUL_3_port) );
  NOR2_X1 U546 ( .A1(n331), .A2(n333), .ZN(Binshift_3_port) );
  INV_X1 U547 ( .A(B[12]), .ZN(n372) );
  INV_X1 U548 ( .A(B[3]), .ZN(n333) );
  NAND4_X1 U549 ( .A1(n359), .A2(n360), .A3(n362), .A4(n363), .ZN(n358) );
  NOR2_X1 U550 ( .A1(n1093), .A2(n359), .ZN(BinLOGIC_19_port) );
  CLKBUF_X1 U551 ( .A(n335), .Z(n1080) );
  AND2_X1 U552 ( .A1(B[15]), .A2(enADDSUB), .ZN(BinADDSUB_15_port) );
  NOR2_X1 U553 ( .A1(n334), .A2(n1091), .ZN(BinLOGIC_2_port) );
  NOR2_X1 U554 ( .A1(n334), .A2(n1097), .ZN(BinMUL_2_port) );
  NOR2_X1 U555 ( .A1(n331), .A2(n334), .ZN(Binshift_2_port) );
  INV_X1 U556 ( .A(B[19]), .ZN(n359) );
  INV_X1 U557 ( .A(B[27]), .ZN(n354) );
  NOR2_X1 U558 ( .A1(n354), .A2(n1086), .ZN(BinADDSUB_27_port) );
  NOR4_X1 U559 ( .A1(n365), .A2(B[10]), .A3(B[12]), .A4(B[11]), .ZN(n341) );
  INV_X1 U560 ( .A(B[28]), .ZN(n356) );
  NOR2_X1 U561 ( .A1(n356), .A2(n1085), .ZN(BinADDSUB_28_port) );
  AND2_X1 U562 ( .A1(B[0]), .A2(enADDSUB), .ZN(BinADDSUB_0_port) );
  NOR2_X1 U564 ( .A1(n360), .A2(n1086), .ZN(BinADDSUB_20_port) );
  AOI22_X1 U570 ( .A1(MULout_25_port), .A2(n1134), .B1(ADDSUBout_25_port), 
        .B2(n1131), .ZN(n107) );
  NOR2_X1 U571 ( .A1(n368), .A2(n1091), .ZN(BinLOGIC_13_port) );
  NOR2_X1 U572 ( .A1(n1098), .A2(n368), .ZN(BinMUL_13_port) );
  AOI22_X1 U573 ( .A1(MULout_29_port), .A2(n1136), .B1(ADDSUBout_29_port), 
        .B2(n1133), .ZN(n309) );
  NOR2_X1 U574 ( .A1(n366), .A2(n1092), .ZN(BinLOGIC_14_port) );
  NOR2_X1 U575 ( .A1(n1097), .A2(n366), .ZN(BinMUL_14_port) );
  NOR2_X1 U576 ( .A1(n350), .A2(n1091), .ZN(BinLOGIC_8_port) );
  NOR2_X1 U577 ( .A1(n1098), .A2(n350), .ZN(BinMUL_8_port) );
  NAND4_X1 U578 ( .A1(n348), .A2(n349), .A3(n350), .A4(n351), .ZN(n347) );
  NOR2_X1 U579 ( .A1(n350), .A2(n1085), .ZN(BinADDSUB_8_port) );
  NOR2_X1 U580 ( .A1(n362), .A2(n1086), .ZN(BinADDSUB_21_port) );
  NOR2_X1 U581 ( .A1(n386), .A2(n1087), .ZN(BinADDSUB_16_port) );
  INV_X1 U582 ( .A(B[16]), .ZN(n386) );
  INV_X1 U583 ( .A(B[10]), .ZN(n375) );
  NOR2_X1 U584 ( .A1(n375), .A2(n1087), .ZN(BinADDSUB_10_port) );
  NOR2_X1 U585 ( .A1(n385), .A2(n1086), .ZN(BinADDSUB_17_port) );
  INV_X1 U586 ( .A(B[17]), .ZN(n385) );
  NOR2_X1 U587 ( .A1(n372), .A2(n1087), .ZN(BinADDSUB_12_port) );
  INV_X1 U588 ( .A(B[15]), .ZN(n367) );
  NOR2_X1 U589 ( .A1(n366), .A2(n1087), .ZN(BinADDSUB_14_port) );
  CLKBUF_X1 U590 ( .A(ADDSUBout_28_port), .Z(n1081) );
  NOR2_X1 U591 ( .A1(n332), .A2(n1085), .ZN(BinADDSUB_4_port) );
  NOR2_X1 U592 ( .A1(n359), .A2(n1086), .ZN(BinADDSUB_19_port) );
  AOI22_X1 U593 ( .A1(MULout_31_port), .A2(n1136), .B1(ADDSUBout_31_port), 
        .B2(n1133), .ZN(n295) );
  INV_X1 U594 ( .A(B[1]), .ZN(n335) );
  NOR2_X1 U595 ( .A1(n348), .A2(n1085), .ZN(BinADDSUB_6_port) );
  INV_X1 U596 ( .A(B[11]), .ZN(n374) );
  NOR2_X1 U597 ( .A1(n367), .A2(n1091), .ZN(BinLOGIC_15_port) );
  NOR2_X1 U598 ( .A1(n1097), .A2(n367), .ZN(BinMUL_15_port) );
  NOR2_X1 U599 ( .A1(n1080), .A2(n1097), .ZN(BinMUL_1_port) );
  NOR2_X1 U600 ( .A1(n1080), .A2(n1092), .ZN(BinLOGIC_1_port) );
  NOR2_X1 U601 ( .A1(n331), .A2(n1080), .ZN(Binshift_1_port) );
  NOR2_X1 U602 ( .A1(n383), .A2(n1086), .ZN(BinADDSUB_23_port) );
  AOI22_X1 U603 ( .A1(MULout_28_port), .A2(n1134), .B1(n1081), .B2(n1131), 
        .ZN(n316) );
  NOR2_X1 U604 ( .A1(n351), .A2(n1085), .ZN(BinADDSUB_9_port) );
  NOR2_X1 U605 ( .A1(n368), .A2(n1087), .ZN(BinADDSUB_13_port) );
  NOR2_X1 U606 ( .A1(n374), .A2(n1087), .ZN(BinADDSUB_11_port) );
  INV_X1 U607 ( .A(B[2]), .ZN(n334) );
  NOR2_X1 U608 ( .A1(n334), .A2(n1085), .ZN(BinADDSUB_2_port) );
  NOR2_X1 U609 ( .A1(n349), .A2(n1085), .ZN(BinADDSUB_7_port) );
  NOR2_X1 U610 ( .A1(n371), .A2(n1085), .ZN(BinADDSUB_5_port) );
  NOR2_X1 U611 ( .A1(n337), .A2(n1091), .ZN(BinLOGIC_0_port) );
  NOR2_X1 U612 ( .A1(n337), .A2(n1097), .ZN(BinMUL_0_port) );
  NOR2_X1 U613 ( .A1(n331), .A2(n337), .ZN(Binshift_0_port) );
  INV_X1 U614 ( .A(B[0]), .ZN(n337) );
  NOR2_X1 U615 ( .A1(n335), .A2(n1086), .ZN(BinADDSUB_1_port) );
  NOR2_X1 U616 ( .A1(n333), .A2(n1085), .ZN(BinADDSUB_3_port) );
  CLKBUF_X1 U617 ( .A(n387), .Z(n1090) );
  CLKBUF_X1 U618 ( .A(n376), .Z(n1096) );
  INV_X1 U619 ( .A(n1079), .ZN(n1113) );
  CLKBUF_X1 U620 ( .A(n1076), .Z(n1127) );
  CLKBUF_X1 U621 ( .A(n1076), .Z(n1128) );
  CLKBUF_X1 U622 ( .A(n1076), .Z(n1129) );
  CLKBUF_X1 U623 ( .A(n1076), .Z(n1130) );
endmodule


module mux21N_N32_9 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   n21, n22, n23, n24;
  assign n21 = S;

  MUX21_470 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n22), .Y(U[0]) );
  MUX21_469 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n24), .Y(U[1]) );
  MUX21_468 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n22), .Y(U[2]) );
  MUX21_467 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n22), .Y(U[3]) );
  MUX21_466 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n22), .Y(U[4]) );
  MUX21_465 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n22), .Y(U[5]) );
  MUX21_464 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n22), .Y(U[6]) );
  MUX21_463 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n22), .Y(U[7]) );
  MUX21_462 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n22), .Y(U[8]) );
  MUX21_461 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n22), .Y(U[9]) );
  MUX21_460 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n22), .Y(U[10]) );
  MUX21_459 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n22), .Y(U[11]) );
  MUX21_458 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n22), .Y(U[12]) );
  MUX21_457 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n23), .Y(U[13]) );
  MUX21_456 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n23), .Y(U[14]) );
  MUX21_455 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n23), .Y(U[15]) );
  MUX21_454 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n23), .Y(U[16]) );
  MUX21_453 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n23), .Y(U[17]) );
  MUX21_452 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n23), .Y(U[18]) );
  MUX21_451 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n23), .Y(U[19]) );
  MUX21_450 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n23), .Y(U[20]) );
  MUX21_449 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n23), .Y(U[21]) );
  MUX21_448 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n23), .Y(U[22]) );
  MUX21_447 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n23), .Y(U[23]) );
  MUX21_446 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n23), .Y(U[24]) );
  MUX21_445 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n24), .Y(U[25]) );
  MUX21_444 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n24), .Y(U[26]) );
  MUX21_443 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n24), .Y(U[27]) );
  MUX21_442 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n24), .Y(U[28]) );
  MUX21_441 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n24), .Y(U[29]) );
  MUX21_440 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n24), .Y(U[30]) );
  MUX21_439 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n24), .Y(U[31]) );
  BUF_X1 U1 ( .A(n21), .Z(n23) );
  BUF_X1 U2 ( .A(n21), .Z(n22) );
  BUF_X1 U3 ( .A(n21), .Z(n24) );
endmodule


module mux41N_Nbit32_0 ( in3, in2, in1, in0, sel, Y );
  input [31:0] in3;
  input [31:0] in2;
  input [31:0] in1;
  input [31:0] in0;
  input [1:0] sel;
  output [31:0] Y;
  wire   \outmux[2][31] , \outmux[2][30] , \outmux[2][29] , \outmux[2][28] ,
         \outmux[2][27] , \outmux[2][26] , \outmux[2][25] , \outmux[2][24] ,
         \outmux[2][23] , \outmux[2][22] , \outmux[2][21] , \outmux[2][20] ,
         \outmux[2][19] , \outmux[2][18] , \outmux[2][17] , \outmux[2][16] ,
         \outmux[2][15] , \outmux[2][14] , \outmux[2][13] , \outmux[2][12] ,
         \outmux[2][11] , \outmux[2][10] , \outmux[2][9] , \outmux[2][8] ,
         \outmux[2][7] , \outmux[2][6] , \outmux[2][5] , \outmux[2][4] ,
         \outmux[2][3] , \outmux[2][2] , \outmux[2][1] , \outmux[2][0] ,
         \outmux[1][31] , \outmux[1][30] , \outmux[1][29] , \outmux[1][28] ,
         \outmux[1][27] , \outmux[1][26] , \outmux[1][25] , \outmux[1][24] ,
         \outmux[1][23] , \outmux[1][22] , \outmux[1][21] , \outmux[1][20] ,
         \outmux[1][19] , \outmux[1][18] , \outmux[1][17] , \outmux[1][16] ,
         \outmux[1][15] , \outmux[1][14] , \outmux[1][13] , \outmux[1][12] ,
         \outmux[1][11] , \outmux[1][10] , \outmux[1][9] , \outmux[1][8] ,
         \outmux[1][7] , \outmux[1][6] , \outmux[1][5] , \outmux[1][4] ,
         \outmux[1][3] , \outmux[1][2] , \outmux[1][1] , \outmux[1][0] ;

  mux21N_N32_6 row1_1 ( .in1(in1), .in0(in0), .S(sel[0]), .U({\outmux[1][31] , 
        \outmux[1][30] , \outmux[1][29] , \outmux[1][28] , \outmux[1][27] , 
        \outmux[1][26] , \outmux[1][25] , \outmux[1][24] , \outmux[1][23] , 
        \outmux[1][22] , \outmux[1][21] , \outmux[1][20] , \outmux[1][19] , 
        \outmux[1][18] , \outmux[1][17] , \outmux[1][16] , \outmux[1][15] , 
        \outmux[1][14] , \outmux[1][13] , \outmux[1][12] , \outmux[1][11] , 
        \outmux[1][10] , \outmux[1][9] , \outmux[1][8] , \outmux[1][7] , 
        \outmux[1][6] , \outmux[1][5] , \outmux[1][4] , \outmux[1][3] , 
        \outmux[1][2] , \outmux[1][1] , \outmux[1][0] }) );
  mux21N_N32_5 row1_2 ( .in1(in3), .in0(in2), .S(sel[0]), .U({\outmux[2][31] , 
        \outmux[2][30] , \outmux[2][29] , \outmux[2][28] , \outmux[2][27] , 
        \outmux[2][26] , \outmux[2][25] , \outmux[2][24] , \outmux[2][23] , 
        \outmux[2][22] , \outmux[2][21] , \outmux[2][20] , \outmux[2][19] , 
        \outmux[2][18] , \outmux[2][17] , \outmux[2][16] , \outmux[2][15] , 
        \outmux[2][14] , \outmux[2][13] , \outmux[2][12] , \outmux[2][11] , 
        \outmux[2][10] , \outmux[2][9] , \outmux[2][8] , \outmux[2][7] , 
        \outmux[2][6] , \outmux[2][5] , \outmux[2][4] , \outmux[2][3] , 
        \outmux[2][2] , \outmux[2][1] , \outmux[2][0] }) );
  mux21N_N32_4 row2_1 ( .in1({\outmux[2][31] , \outmux[2][30] , 
        \outmux[2][29] , \outmux[2][28] , \outmux[2][27] , \outmux[2][26] , 
        \outmux[2][25] , \outmux[2][24] , \outmux[2][23] , \outmux[2][22] , 
        \outmux[2][21] , \outmux[2][20] , \outmux[2][19] , \outmux[2][18] , 
        \outmux[2][17] , \outmux[2][16] , \outmux[2][15] , \outmux[2][14] , 
        \outmux[2][13] , \outmux[2][12] , \outmux[2][11] , \outmux[2][10] , 
        \outmux[2][9] , \outmux[2][8] , \outmux[2][7] , \outmux[2][6] , 
        \outmux[2][5] , \outmux[2][4] , \outmux[2][3] , \outmux[2][2] , 
        \outmux[2][1] , \outmux[2][0] }), .in0({\outmux[1][31] , 
        \outmux[1][30] , \outmux[1][29] , \outmux[1][28] , \outmux[1][27] , 
        \outmux[1][26] , \outmux[1][25] , \outmux[1][24] , \outmux[1][23] , 
        \outmux[1][22] , \outmux[1][21] , \outmux[1][20] , \outmux[1][19] , 
        \outmux[1][18] , \outmux[1][17] , \outmux[1][16] , \outmux[1][15] , 
        \outmux[1][14] , \outmux[1][13] , \outmux[1][12] , \outmux[1][11] , 
        \outmux[1][10] , \outmux[1][9] , \outmux[1][8] , \outmux[1][7] , 
        \outmux[1][6] , \outmux[1][5] , \outmux[1][4] , \outmux[1][3] , 
        \outmux[1][2] , \outmux[1][1] , \outmux[1][0] }), .S(sel[1]), .U(Y) );
endmodule


module mux21N_N32_10 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   n14, n15, n16, n17;
  tri   net389393;
  assign net389393 = S;

  MUX21_502 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n14), .Y(U[0]) );
  MUX21_501 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n17), .Y(U[1]) );
  MUX21_500 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n16), .Y(U[2]) );
  MUX21_499 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n14), .Y(U[3]) );
  MUX21_498 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n17), .Y(U[4]) );
  MUX21_497 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n16), .Y(U[5]) );
  MUX21_496 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n15), .Y(U[6]) );
  MUX21_495 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n17), .Y(U[7]) );
  MUX21_494 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n15), .Y(U[8]) );
  MUX21_493 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n17), .Y(U[9]) );
  MUX21_492 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n16), .Y(U[10]) );
  MUX21_491 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n15), .Y(U[11]) );
  MUX21_490 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n16), .Y(U[12]) );
  MUX21_489 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n16), .Y(U[13]) );
  MUX21_488 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n17), .Y(U[14]) );
  MUX21_487 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n15), .Y(U[15]) );
  MUX21_486 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n15), .Y(U[16]) );
  MUX21_485 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n15), .Y(U[17]) );
  MUX21_484 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n16), .Y(U[18]) );
  MUX21_483 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n16), .Y(U[19]) );
  MUX21_482 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n15), .Y(U[20]) );
  MUX21_481 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n17), .Y(U[21]) );
  MUX21_480 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n17), .Y(U[22]) );
  MUX21_479 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n17), .Y(U[23]) );
  MUX21_478 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n16), .Y(U[24]) );
  MUX21_477 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n17), .Y(U[25]) );
  MUX21_476 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n15), .Y(U[26]) );
  MUX21_475 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n15), .Y(U[27]) );
  MUX21_474 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n16), .Y(U[28]) );
  MUX21_473 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n17), .Y(U[29]) );
  MUX21_472 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n15), .Y(U[30]) );
  MUX21_471 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n16), .Y(U[31]) );
  BUF_X2 U1 ( .A(net389393), .Z(n16) );
  BUF_X2 U2 ( .A(net389393), .Z(n15) );
  BUF_X2 U3 ( .A(net389393), .Z(n17) );
  CLKBUF_X1 U4 ( .A(net389393), .Z(n14) );
endmodule


module FD_EN_435 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module RegEn_Nbit32_5 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;


  FD_EN_170 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_169 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_168 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_167 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_166 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
  FD_EN_165 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[5]) );
  FD_EN_164 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[6]) );
  FD_EN_163 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[7]) );
  FD_EN_162 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[8]) );
  FD_EN_161 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[9]) );
  FD_EN_160 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[10])
         );
  FD_EN_159 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[11])
         );
  FD_EN_158 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[12])
         );
  FD_EN_157 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[13])
         );
  FD_EN_156 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[14])
         );
  FD_EN_155 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[15])
         );
  FD_EN_154 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[16])
         );
  FD_EN_153 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[17])
         );
  FD_EN_152 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[18])
         );
  FD_EN_151 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[19])
         );
  FD_EN_150 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[20])
         );
  FD_EN_149 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[21])
         );
  FD_EN_148 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[22])
         );
  FD_EN_147 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[23])
         );
  FD_EN_146 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[24])
         );
  FD_EN_145 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[25])
         );
  FD_EN_144 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[26])
         );
  FD_EN_143 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[27])
         );
  FD_EN_142 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[28])
         );
  FD_EN_141 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[29])
         );
  FD_EN_140 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[30])
         );
  FD_EN_139 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[31])
         );
endmodule


module RegEn_Nbit32_6 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;


  FD_EN_202 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_201 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_200 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_199 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_198 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
  FD_EN_197 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[5]) );
  FD_EN_196 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[6]) );
  FD_EN_195 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[7]) );
  FD_EN_194 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[8]) );
  FD_EN_193 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[9]) );
  FD_EN_192 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[10])
         );
  FD_EN_191 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[11])
         );
  FD_EN_190 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[12])
         );
  FD_EN_189 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[13])
         );
  FD_EN_188 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[14])
         );
  FD_EN_187 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[15])
         );
  FD_EN_186 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[16])
         );
  FD_EN_185 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[17])
         );
  FD_EN_184 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[18])
         );
  FD_EN_183 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[19])
         );
  FD_EN_182 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[20])
         );
  FD_EN_181 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[21])
         );
  FD_EN_180 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[22])
         );
  FD_EN_179 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[23])
         );
  FD_EN_178 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[24])
         );
  FD_EN_177 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[25])
         );
  FD_EN_176 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[26])
         );
  FD_EN_175 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[27])
         );
  FD_EN_174 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[28])
         );
  FD_EN_173 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[29])
         );
  FD_EN_172 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[30])
         );
  FD_EN_171 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[31])
         );
endmodule


module RegEn_Nbit5_0 ( A, Clk, Reset, EN, U );
  input [4:0] A;
  output [4:0] U;
  input Clk, Reset, EN;


  FD_EN_207 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_206 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_205 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_204 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_203 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
endmodule


module RegEn_Nbit32_7 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;


  FD_EN_239 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_238 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_237 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_236 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_235 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
  FD_EN_234 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[5]) );
  FD_EN_233 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[6]) );
  FD_EN_232 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[7]) );
  FD_EN_231 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[8]) );
  FD_EN_230 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[9]) );
  FD_EN_229 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[10])
         );
  FD_EN_228 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[11])
         );
  FD_EN_227 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[12])
         );
  FD_EN_226 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[13])
         );
  FD_EN_225 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[14])
         );
  FD_EN_224 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[15])
         );
  FD_EN_223 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[16])
         );
  FD_EN_222 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[17])
         );
  FD_EN_221 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[18])
         );
  FD_EN_220 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[19])
         );
  FD_EN_219 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[20])
         );
  FD_EN_218 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[21])
         );
  FD_EN_217 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[22])
         );
  FD_EN_216 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[23])
         );
  FD_EN_215 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[24])
         );
  FD_EN_214 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[25])
         );
  FD_EN_213 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[26])
         );
  FD_EN_212 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[27])
         );
  FD_EN_211 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[28])
         );
  FD_EN_210 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[29])
         );
  FD_EN_209 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[30])
         );
  FD_EN_208 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[31])
         );
endmodule


module RegEn_Nbit32_8 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;

  tri   [31:0] A;

  FD_EN_271 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_270 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_269 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_268 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_267 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
  FD_EN_266 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[5]) );
  FD_EN_265 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[6]) );
  FD_EN_264 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[7]) );
  FD_EN_263 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[8]) );
  FD_EN_262 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[9]) );
  FD_EN_261 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[10])
         );
  FD_EN_260 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[11])
         );
  FD_EN_259 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[12])
         );
  FD_EN_258 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[13])
         );
  FD_EN_257 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[14])
         );
  FD_EN_256 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[15])
         );
  FD_EN_255 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[16])
         );
  FD_EN_254 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[17])
         );
  FD_EN_253 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[18])
         );
  FD_EN_252 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[19])
         );
  FD_EN_251 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[20])
         );
  FD_EN_250 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[21])
         );
  FD_EN_249 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[22])
         );
  FD_EN_248 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[23])
         );
  FD_EN_247 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[24])
         );
  FD_EN_246 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[25])
         );
  FD_EN_245 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[26])
         );
  FD_EN_244 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[27])
         );
  FD_EN_243 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[28])
         );
  FD_EN_242 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[29])
         );
  FD_EN_241 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[30])
         );
  FD_EN_240 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[31])
         );
endmodule


module RegEn_Nbit32_9 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;

  tri   [31:0] A;

  FD_EN_303 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_302 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_301 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_300 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_299 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
  FD_EN_298 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[5]) );
  FD_EN_297 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[6]) );
  FD_EN_296 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[7]) );
  FD_EN_295 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[8]) );
  FD_EN_294 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[9]) );
  FD_EN_293 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[10])
         );
  FD_EN_292 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[11])
         );
  FD_EN_291 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[12])
         );
  FD_EN_290 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[13])
         );
  FD_EN_289 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[14])
         );
  FD_EN_288 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[15])
         );
  FD_EN_287 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[16])
         );
  FD_EN_286 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[17])
         );
  FD_EN_285 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[18])
         );
  FD_EN_284 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[19])
         );
  FD_EN_283 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[20])
         );
  FD_EN_282 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[21])
         );
  FD_EN_281 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[22])
         );
  FD_EN_280 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[23])
         );
  FD_EN_279 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[24])
         );
  FD_EN_278 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[25])
         );
  FD_EN_277 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[26])
         );
  FD_EN_276 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[27])
         );
  FD_EN_275 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[28])
         );
  FD_EN_274 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[29])
         );
  FD_EN_273 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[30])
         );
  FD_EN_272 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[31])
         );
endmodule


module FD_EN_436 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module mux21N_N32_11 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   n21, n22, n23, n24;
  assign n21 = S;

  MUX21_534 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n22), .Y(U[0]) );
  MUX21_533 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n22), .Y(U[1]) );
  MUX21_532 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n22), .Y(U[2]) );
  MUX21_531 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n22), .Y(U[3]) );
  MUX21_530 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n22), .Y(U[4]) );
  MUX21_529 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n22), .Y(U[5]) );
  MUX21_528 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n22), .Y(U[6]) );
  MUX21_527 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n22), .Y(U[7]) );
  MUX21_526 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n22), .Y(U[8]) );
  MUX21_525 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n22), .Y(U[9]) );
  MUX21_524 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n22), .Y(U[10]) );
  MUX21_523 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n22), .Y(U[11]) );
  MUX21_522 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n23), .Y(U[12]) );
  MUX21_521 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n23), .Y(U[13]) );
  MUX21_520 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n23), .Y(U[14]) );
  MUX21_519 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n23), .Y(U[15]) );
  MUX21_518 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n23), .Y(U[16]) );
  MUX21_517 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n23), .Y(U[17]) );
  MUX21_516 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n23), .Y(U[18]) );
  MUX21_515 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n23), .Y(U[19]) );
  MUX21_514 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n23), .Y(U[20]) );
  MUX21_513 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n23), .Y(U[21]) );
  MUX21_512 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n23), .Y(U[22]) );
  MUX21_511 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n23), .Y(U[23]) );
  MUX21_510 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n24), .Y(U[24]) );
  MUX21_509 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n24), .Y(U[25]) );
  MUX21_508 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n24), .Y(U[26]) );
  MUX21_507 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n24), .Y(U[27]) );
  MUX21_506 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n24), .Y(U[28]) );
  MUX21_505 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n24), .Y(U[29]) );
  MUX21_504 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n24), .Y(U[30]) );
  MUX21_503 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n24), .Y(U[31]) );
  BUF_X1 U1 ( .A(n21), .Z(n23) );
  BUF_X1 U2 ( .A(n21), .Z(n22) );
  BUF_X1 U3 ( .A(n21), .Z(n24) );
endmodule


module zerotest_Nbit32 ( A, zero );
  input [31:0] A;
  output zero;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  tri   [31:0] A;

  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(zero) );
  NOR4_X1 U2 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n6) );
  NOR4_X1 U3 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n10) );
  NAND4_X1 U4 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NOR4_X1 U5 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n3) );
  NOR4_X1 U6 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n4) );
  NOR4_X1 U7 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n5) );
  NAND4_X1 U8 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
  NOR4_X1 U9 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n7) );
  NOR4_X1 U10 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n8) );
  NOR4_X1 U11 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n9) );
endmodule


module mux21N_N32_12 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   n21, n22, n23, n24;
  tri   [31:0] in1;
  assign n21 = S;

  MUX21_566 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n22), .Y(U[0]) );
  MUX21_565 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n22), .Y(U[1]) );
  MUX21_564 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n22), .Y(U[2]) );
  MUX21_563 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n22), .Y(U[3]) );
  MUX21_562 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n22), .Y(U[4]) );
  MUX21_561 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n22), .Y(U[5]) );
  MUX21_560 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n22), .Y(U[6]) );
  MUX21_559 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n22), .Y(U[7]) );
  MUX21_558 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n22), .Y(U[8]) );
  MUX21_557 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n22), .Y(U[9]) );
  MUX21_556 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n22), .Y(U[10]) );
  MUX21_555 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n22), .Y(U[11]) );
  MUX21_554 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n23), .Y(U[12]) );
  MUX21_553 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n23), .Y(U[13]) );
  MUX21_552 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n23), .Y(U[14]) );
  MUX21_551 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n23), .Y(U[15]) );
  MUX21_550 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n23), .Y(U[16]) );
  MUX21_549 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n23), .Y(U[17]) );
  MUX21_548 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n23), .Y(U[18]) );
  MUX21_547 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n23), .Y(U[19]) );
  MUX21_546 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n23), .Y(U[20]) );
  MUX21_545 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n23), .Y(U[21]) );
  MUX21_544 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n23), .Y(U[22]) );
  MUX21_543 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n23), .Y(U[23]) );
  MUX21_542 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n24), .Y(U[24]) );
  MUX21_541 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n24), .Y(U[25]) );
  MUX21_540 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n24), .Y(U[26]) );
  MUX21_539 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n24), .Y(U[27]) );
  MUX21_538 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n24), .Y(U[28]) );
  MUX21_537 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n24), .Y(U[29]) );
  MUX21_536 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n24), .Y(U[30]) );
  MUX21_535 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n24), .Y(U[31]) );
  BUF_X1 U1 ( .A(n21), .Z(n23) );
  BUF_X1 U2 ( .A(n21), .Z(n22) );
  BUF_X1 U3 ( .A(n21), .Z(n24) );
endmodule


module AddSubN_Nbit32_2 ( A, B, addnsub, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input addnsub;
  output Cout;

  wire   [31:0] addendB;
  wire   [7:0] Carry;

  SparseTreeCarryGenN_Nbit32_2 STCG ( .A(A), .B(addendB), .Cin(addnsub), 
        .Cout({Cout, Carry}) );
  CarrySumN_Nbit32_2 CSN ( .A(A), .B(addendB), .Ci(Carry), .S(S) );
  XOR2_X1 U1 ( .A(addnsub), .B(B[9]), .Z(addendB[9]) );
  XOR2_X1 U2 ( .A(addnsub), .B(B[8]), .Z(addendB[8]) );
  XOR2_X1 U3 ( .A(addnsub), .B(B[7]), .Z(addendB[7]) );
  XOR2_X1 U4 ( .A(addnsub), .B(B[6]), .Z(addendB[6]) );
  XOR2_X1 U5 ( .A(addnsub), .B(B[5]), .Z(addendB[5]) );
  XOR2_X1 U6 ( .A(addnsub), .B(B[4]), .Z(addendB[4]) );
  XOR2_X1 U7 ( .A(addnsub), .B(B[3]), .Z(addendB[3]) );
  XOR2_X1 U8 ( .A(addnsub), .B(B[31]), .Z(addendB[31]) );
  XOR2_X1 U9 ( .A(addnsub), .B(B[30]), .Z(addendB[30]) );
  XOR2_X1 U10 ( .A(addnsub), .B(B[2]), .Z(addendB[2]) );
  XOR2_X1 U11 ( .A(addnsub), .B(B[29]), .Z(addendB[29]) );
  XOR2_X1 U12 ( .A(addnsub), .B(B[28]), .Z(addendB[28]) );
  XOR2_X1 U13 ( .A(addnsub), .B(B[27]), .Z(addendB[27]) );
  XOR2_X1 U14 ( .A(addnsub), .B(B[26]), .Z(addendB[26]) );
  XOR2_X1 U15 ( .A(addnsub), .B(B[25]), .Z(addendB[25]) );
  XOR2_X1 U16 ( .A(addnsub), .B(B[24]), .Z(addendB[24]) );
  XOR2_X1 U17 ( .A(addnsub), .B(B[23]), .Z(addendB[23]) );
  XOR2_X1 U18 ( .A(addnsub), .B(B[22]), .Z(addendB[22]) );
  XOR2_X1 U19 ( .A(addnsub), .B(B[21]), .Z(addendB[21]) );
  XOR2_X1 U20 ( .A(addnsub), .B(B[20]), .Z(addendB[20]) );
  XOR2_X1 U21 ( .A(addnsub), .B(B[1]), .Z(addendB[1]) );
  XOR2_X1 U22 ( .A(addnsub), .B(B[19]), .Z(addendB[19]) );
  XOR2_X1 U23 ( .A(addnsub), .B(B[18]), .Z(addendB[18]) );
  XOR2_X1 U24 ( .A(addnsub), .B(B[17]), .Z(addendB[17]) );
  XOR2_X1 U25 ( .A(addnsub), .B(B[16]), .Z(addendB[16]) );
  XOR2_X1 U26 ( .A(addnsub), .B(B[15]), .Z(addendB[15]) );
  XOR2_X1 U27 ( .A(addnsub), .B(B[14]), .Z(addendB[14]) );
  XOR2_X1 U28 ( .A(addnsub), .B(B[13]), .Z(addendB[13]) );
  XOR2_X1 U29 ( .A(addnsub), .B(B[12]), .Z(addendB[12]) );
  XOR2_X1 U30 ( .A(addnsub), .B(B[11]), .Z(addendB[11]) );
  XOR2_X1 U31 ( .A(addnsub), .B(B[10]), .Z(addendB[10]) );
  XOR2_X1 U32 ( .A(addnsub), .B(B[0]), .Z(addendB[0]) );
endmodule


module signExtension_Nbitin26_Nbitout32 ( A, Aextended );
  input [25:0] A;
  output [31:0] Aextended;

  assign Aextended[31] = A[25];
  assign Aextended[30] = A[25];
  assign Aextended[29] = A[25];
  assign Aextended[28] = A[25];
  assign Aextended[27] = A[25];
  assign Aextended[26] = A[25];
  assign Aextended[25] = A[25];
  assign Aextended[24] = A[24];
  assign Aextended[23] = A[23];
  assign Aextended[22] = A[22];
  assign Aextended[21] = A[21];
  assign Aextended[20] = A[20];
  assign Aextended[19] = A[19];
  assign Aextended[18] = A[18];
  assign Aextended[17] = A[17];
  assign Aextended[16] = A[16];
  assign Aextended[15] = A[15];
  assign Aextended[14] = A[14];
  assign Aextended[13] = A[13];
  assign Aextended[12] = A[12];
  assign Aextended[11] = A[11];
  assign Aextended[10] = A[10];
  assign Aextended[9] = A[9];
  assign Aextended[8] = A[8];
  assign Aextended[7] = A[7];
  assign Aextended[6] = A[6];
  assign Aextended[5] = A[5];
  assign Aextended[4] = A[4];
  assign Aextended[3] = A[3];
  assign Aextended[2] = A[2];
  assign Aextended[1] = A[1];
  assign Aextended[0] = A[0];

endmodule


module signExtension_Nbitin16_Nbitout32_1 ( A, Aextended );
  input [15:0] A;
  output [31:0] Aextended;

  assign Aextended[31] = A[15];
  assign Aextended[30] = A[15];
  assign Aextended[29] = A[15];
  assign Aextended[28] = A[15];
  assign Aextended[27] = A[15];
  assign Aextended[26] = A[15];
  assign Aextended[25] = A[15];
  assign Aextended[24] = A[15];
  assign Aextended[23] = A[15];
  assign Aextended[22] = A[15];
  assign Aextended[21] = A[15];
  assign Aextended[20] = A[15];
  assign Aextended[19] = A[15];
  assign Aextended[18] = A[15];
  assign Aextended[17] = A[15];
  assign Aextended[16] = A[15];
  assign Aextended[15] = A[15];
  assign Aextended[14] = A[14];
  assign Aextended[13] = A[13];
  assign Aextended[12] = A[12];
  assign Aextended[11] = A[11];
  assign Aextended[10] = A[10];
  assign Aextended[9] = A[9];
  assign Aextended[8] = A[8];
  assign Aextended[7] = A[7];
  assign Aextended[6] = A[6];
  assign Aextended[5] = A[5];
  assign Aextended[4] = A[4];
  assign Aextended[3] = A[3];
  assign Aextended[2] = A[2];
  assign Aextended[1] = A[1];
  assign Aextended[0] = A[0];

endmodule


module signExtension_Nbitin16_Nbitout32_0 ( A, Aextended );
  input [15:0] A;
  output [31:0] Aextended;

  assign Aextended[31] = A[15];
  assign Aextended[30] = A[15];
  assign Aextended[29] = A[15];
  assign Aextended[28] = A[15];
  assign Aextended[27] = A[15];
  assign Aextended[26] = A[15];
  assign Aextended[25] = A[15];
  assign Aextended[24] = A[15];
  assign Aextended[23] = A[15];
  assign Aextended[22] = A[15];
  assign Aextended[21] = A[15];
  assign Aextended[20] = A[15];
  assign Aextended[19] = A[15];
  assign Aextended[18] = A[15];
  assign Aextended[17] = A[15];
  assign Aextended[16] = A[15];
  assign Aextended[15] = A[15];
  assign Aextended[14] = A[14];
  assign Aextended[13] = A[13];
  assign Aextended[12] = A[12];
  assign Aextended[11] = A[11];
  assign Aextended[10] = A[10];
  assign Aextended[9] = A[9];
  assign Aextended[8] = A[8];
  assign Aextended[7] = A[7];
  assign Aextended[6] = A[6];
  assign Aextended[5] = A[5];
  assign Aextended[4] = A[4];
  assign Aextended[3] = A[3];
  assign Aextended[2] = A[2];
  assign Aextended[1] = A[1];
  assign Aextended[0] = A[0];

endmodule


module register_file_Nbit32 ( CLK, RESET, ENABLE, RD1, RD2, WR, ADD_WR, 
        ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5457, n5459, n5461, n5463, n5465, n5467, n5469,
         n5471, n5472, n5473, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4977, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n18773, n18776, n1078, n1079, n1080, n1083,
         n1085, n1087, n1089, n1091, n1093, n1095, n1097, n1099, n1101, n1103,
         n1105, n1107, n1109, n1111, n1113, n1115, n1117, n1119, n1121, n1123,
         n1125, n1127, n1129, n1131, n1133, n1135, n1137, n1139, n1141, n1143,
         n1145, n1146, n1148, n1149, n1150, n1151, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1225, n1226, n1227, n1260, n1263, n1295, n1297,
         n1298, n1301, n1335, n1367, n1368, n1371, n1403, n1405, n1437, n1439,
         n1440, n1441, n1443, n1444, n1446, n1447, n1450, n1484, n1517, n1520,
         n1554, n1586, n1589, n1623, n1655, n1657, n1658, n1661, n1695, n1727,
         n1730, n1764, n1796, n1799, n1833, n1834, n1835, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1858, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1870, n1871, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1889, n1890, n1891, n1892, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1908, n1909, n1912, n1913, n1914, n1915, n1917, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1933,
         n1934, n1937, n1938, n1939, n1940, n1942, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1958, n1959,
         n1962, n1963, n1964, n1965, n1967, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1983, n1984, n1987,
         n1988, n1989, n1990, n1992, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2008, n2009, n2012, n2013,
         n2014, n2015, n2017, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2033, n2034, n2037, n2038, n2039,
         n2040, n2042, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2058, n2059, n2062, n2063, n2064, n2065,
         n2067, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2083, n2084, n2087, n2088, n2089, n2090, n2092,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2108, n2109, n2112, n2113, n2114, n2115, n2117, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2133, n2134, n2137, n2138, n2139, n2140, n2142, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2158, n2159, n2162, n2163, n2164, n2165, n2167, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2183,
         n2184, n2187, n2188, n2189, n2190, n2192, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2208, n2209,
         n2212, n2213, n2214, n2215, n2217, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2233, n2234, n2237,
         n2238, n2239, n2240, n2242, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2258, n2259, n2262, n2263,
         n2264, n2265, n2267, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2283, n2284, n2287, n2288, n2289,
         n2290, n2292, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2308, n2309, n2312, n2313, n2314, n2315,
         n2317, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2333, n2334, n2337, n2338, n2339, n2340, n2342,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2358, n2359, n2362, n2363, n2364, n2365, n2367, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2383, n2384, n2387, n2388, n2389, n2390, n2392, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2408, n2409, n2412, n2413, n2414, n2415, n2417, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2433,
         n2434, n2437, n2438, n2439, n2440, n2442, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2458, n2459,
         n2462, n2463, n2464, n2465, n2467, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2483, n2484, n2487,
         n2488, n2489, n2490, n2492, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2508, n2509, n2512, n2513,
         n2514, n2515, n2517, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2533, n2534, n2537, n2538, n2539,
         n2540, n2542, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2558, n2559, n2562, n2563, n2564, n2565,
         n2567, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2583, n2584, n2587, n2588, n2589, n2590, n2592,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2608, n2609, n2612, n2613, n2614, n2615, n2617, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2633, n2634, n2637, n2638, n2639, n2640, n2642, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2673, n2674, n2675, n2676, n2677,
         n2678, n2680, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2723, n2724, n2725, n2726, n2727, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2765, n2767, n2768, n2769, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2787,
         n2789, n2790, n2791, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2809, n2811,
         n2812, n2813, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2831, n2833, n2834,
         n2835, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2853, n2855, n2856, n2857,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2875, n2877, n2878, n2879, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2897, n2899, n2900, n2901, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2919, n2921, n2922, n2923, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2941, n2943, n2944, n2945, n2947, n2948, n2949, n2950,
         n2951, n2952, n3081, n3082, n4395, n4460, n4461, n4462, n4463, n4464,
         n4465, n4467, n4469, n4470, n4471, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4489, n4491, n4492, n4493, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4511,
         n4513, n4514, n4515, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4533, n4535,
         n4536, n4537, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4555, n4557, n4558,
         n4559, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4577, n4579, n4580, n4581,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4599, n4601, n4602, n4603, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4621, n4623, n4624, n4625, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4643, n4645, n4646, n4647, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4665, n4667, n4668, n4669, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4687, n4689, n4690, n4691, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4709, n4711, n4712, n4713, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4731,
         n4733, n4734, n4735, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4753, n4755,
         n4756, n4757, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4775, n4777, n4778,
         n4875, n4877, n4878, n4879, n4880, n4881, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4907, n4909, n4910, n4911,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4942, n4944, n4945, n4946, n4948,
         n4949, n4950, n4951, n4976, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5313, n5315, n5316, n5317, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5631, n5633, n5634, n5635, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5653, n5655, n5656, n5657, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5675, n5677, n5678, n5679, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5706,
         n5707, n5708, n5710, n5711, n5712, n5713, n5714, n5715, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758;
  tri   RD1;
  tri   RD2;
  tri   WR;
  tri   [31:0] OUT1;
  tri   [31:0] OUT2;

  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(n4394), .CK(CLK), .RN(n20732), .Q(n5620), 
        .QN(n19026) );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(n4393), .CK(CLK), .RN(n20718), .Q(n5619), 
        .QN(n19032) );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(n4392), .CK(CLK), .RN(n20696), .Q(n5618), 
        .QN(n19040) );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(n4391), .CK(CLK), .RN(n20740), .Q(n5617), 
        .QN(n19025) );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(n4390), .CK(CLK), .RN(n20705), .Q(n5616), 
        .QN(n19031) );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(n4389), .CK(CLK), .RN(n20692), .Q(n5615), 
        .QN(n19039) );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(n4388), .CK(CLK), .RN(n20708), .Q(n5614), 
        .QN(n19024) );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(n4387), .CK(CLK), .RN(n20699), .Q(n5613), 
        .QN(n19023) );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(n4386), .CK(CLK), .RN(n20741), .Q(n5612), 
        .QN(n19042) );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(n4385), .CK(CLK), .RN(n20700), .Q(n5611), 
        .QN(n19022) );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(n4384), .CK(CLK), .RN(n20709), .Q(n5630), 
        .QN(n19021) );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(n4383), .CK(CLK), .RN(n20719), .Q(n5629), 
        .QN(n19038) );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(n4382), .CK(CLK), .RN(n20727), .Q(n5610), 
        .QN(n19020) );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(n4381), .CK(CLK), .RN(n20739), .Q(n5609), 
        .QN(n19019) );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(n4380), .CK(CLK), .RN(n20697), .Q(n5608), 
        .QN(n19037) );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(n4379), .CK(CLK), .RN(n20735), .Q(n5607), 
        .QN(n19030) );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(n4378), .CK(CLK), .RN(n20694), .Q(n5606), 
        .QN(n19018) );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(n4377), .CK(CLK), .RN(n20701), .Q(n5605), 
        .QN(n19036) );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(n4376), .CK(CLK), .RN(n20730), .Q(n5604), 
        .QN(n19017) );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(n4375), .CK(CLK), .RN(n20702), .Q(n5603), 
        .QN(n19029) );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(n4374), .CK(CLK), .RN(n20692), .Q(n5415), 
        .QN(n19035) );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(n4373), .CK(CLK), .RN(n20727), .Q(n5414), 
        .QN(n19016) );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(n4372), .CK(CLK), .RN(n20710), .Q(n5413), 
        .QN(n19028) );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(n4371), .CK(CLK), .RN(n20733), .Q(n5412), 
        .QN(n19034) );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(n4370), .CK(CLK), .RN(n20723), .Q(n5411), 
        .QN(n19015) );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(n4369), .CK(CLK), .RN(n20711), .Q(n5410), 
        .QN(n19014) );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(n4368), .CK(CLK), .RN(n20696), .Q(n5409), 
        .QN(n19041) );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(n4367), .CK(CLK), .RN(n20703), .Q(n5408), 
        .QN(n19013) );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(n4366), .CK(CLK), .RN(n20720), .Q(n5407), 
        .QN(n19012) );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(n4365), .CK(CLK), .RN(n20712), .Q(n5406), 
        .QN(n19033) );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(n4364), .CK(CLK), .RN(n20694), .Q(n5405), 
        .QN(n19027) );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(n4363), .CK(CLK), .RN(n20737), .Q(n5404), 
        .QN(n19011) );
  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(n4362), .CK(CLK), .RN(n20720), .Q(n19490), .QN(n4874) );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(n4361), .CK(CLK), .RN(n20715), .Q(n19489), .QN(n4873) );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(n4360), .CK(CLK), .RN(n20710), .Q(n19488), .QN(n4872) );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(n4359), .CK(CLK), .RN(n20744), .Q(n19487), .QN(n4871) );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(n4358), .CK(CLK), .RN(n20740), .Q(n19486), .QN(n4870) );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(n4357), .CK(CLK), .RN(n20727), .Q(n19485), .QN(n4869) );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(n4356), .CK(CLK), .RN(n20699), .Q(n19484), .QN(n4868) );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(n4355), .CK(CLK), .RN(n20698), .Q(n19483), .QN(n4867) );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(n4354), .CK(CLK), .RN(n20718), .Q(n19482), .QN(n4866) );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(n4353), .CK(CLK), .RN(n20705), .Q(n19481), .QN(n4865) );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(n4352), .CK(CLK), .RN(n20696), .Q(n19480), .QN(n4864) );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(n4351), .CK(CLK), .RN(n20697), .Q(n19479), .QN(n4863) );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(n4350), .CK(CLK), .RN(n20717), .Q(n19478), .QN(n4862) );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(n4349), .CK(CLK), .RN(n20697), .Q(n19477), .QN(n4861) );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(n4348), .CK(CLK), .RN(n20703), .Q(n19476), .QN(n4860) );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(n4347), .CK(CLK), .RN(n20718), .Q(n19475), .QN(n4859) );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(n4346), .CK(CLK), .RN(n20694), .Q(n19474), .QN(n4858) );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(n4345), .CK(CLK), .RN(n20700), .Q(n19473), .QN(n4857) );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(n4344), .CK(CLK), .RN(n20701), .Q(n19472), .QN(n4856) );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(n4343), .CK(CLK), .RN(n20716), .Q(n19471), .QN(n4855) );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(n4342), .CK(CLK), .RN(n20727), .Q(n19470), .QN(n4854) );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(n4341), .CK(CLK), .RN(n20741), .Q(n19469), .QN(n4853) );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(n4340), .CK(CLK), .RN(n20741), .Q(n19468), 
        .QN(n4852) );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(n4339), .CK(CLK), .RN(n20691), .Q(n19467), 
        .QN(n4851) );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(n4338), .CK(CLK), .RN(n20742), .Q(n19466), 
        .QN(n4850) );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(n4337), .CK(CLK), .RN(n20745), .Q(n19465), 
        .QN(n4849) );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(n4336), .CK(CLK), .RN(n20725), .Q(n19464), 
        .QN(n4848) );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(n4335), .CK(CLK), .RN(n20714), .Q(n19463), 
        .QN(n4847) );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(n4334), .CK(CLK), .RN(n20734), .Q(n19462), 
        .QN(n4846) );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(n4333), .CK(CLK), .RN(n20709), .Q(n19461), 
        .QN(n4845) );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(n4332), .CK(CLK), .RN(n20704), .Q(n19460), 
        .QN(n4844) );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(n4331), .CK(CLK), .RN(n20719), .Q(n19459), 
        .QN(n4843) );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(n4330), .CK(CLK), .RN(n20705), .Q(n5403), 
        .QN(n19234) );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(n4329), .CK(CLK), .RN(n20691), .Q(n5402), 
        .QN(n19233) );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(n4328), .CK(CLK), .RN(n20697), .Q(n5401), 
        .QN(n19232) );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(n4327), .CK(CLK), .RN(n20744), .Q(n5400), 
        .QN(n19231) );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(n4326), .CK(CLK), .RN(n20710), .Q(n5399), 
        .QN(n19230) );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(n4325), .CK(CLK), .RN(n20736), .Q(n5398), 
        .QN(n19229) );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(n4324), .CK(CLK), .RN(n20692), .Q(n5397), 
        .QN(n19228) );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(n4323), .CK(CLK), .RN(n20698), .Q(n5396), 
        .QN(n19227) );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(n4322), .CK(CLK), .RN(n20734), .Q(n5395), 
        .QN(n19226) );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(n4321), .CK(CLK), .RN(n20731), .Q(n5394), 
        .QN(n19225) );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(n4320), .CK(CLK), .RN(n20692), .Q(n5393), 
        .QN(n19224) );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(n4319), .CK(CLK), .RN(n20719), .Q(n5392), 
        .QN(n19223) );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(n4318), .CK(CLK), .RN(n20717), .Q(n5391), 
        .QN(n19222) );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(n4317), .CK(CLK), .RN(n20724), .Q(n5390), 
        .QN(n19221) );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(n4316), .CK(CLK), .RN(n20711), .Q(n5389), 
        .QN(n19220) );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(n4315), .CK(CLK), .RN(n20704), .Q(n5388), 
        .QN(n19219) );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(n4314), .CK(CLK), .RN(n20694), .Q(n5387), 
        .QN(n19218) );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(n4313), .CK(CLK), .RN(n20727), .Q(n5386), 
        .QN(n19217) );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(n4312), .CK(CLK), .RN(n20699), .Q(n5385), 
        .QN(n19216) );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(n4311), .CK(CLK), .RN(n20716), .Q(n5384), 
        .QN(n19215) );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(n4310), .CK(CLK), .RN(n20741), .Q(n5301), 
        .QN(n19214) );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(n4309), .CK(CLK), .RN(n20692), .Q(n5300), 
        .QN(n19213) );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(n4308), .CK(CLK), .RN(n20710), .Q(n5299), 
        .QN(n19212) );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(n4307), .CK(CLK), .RN(n20691), .Q(n5298), 
        .QN(n19211) );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(n4306), .CK(CLK), .RN(n20742), .Q(n5297), 
        .QN(n19210) );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(n4305), .CK(CLK), .RN(n20708), .Q(n5296), 
        .QN(n19209) );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(n4304), .CK(CLK), .RN(n20725), .Q(n5295), 
        .QN(n19208) );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(n4303), .CK(CLK), .RN(n20712), .Q(n5294), 
        .QN(n19207) );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(n4302), .CK(CLK), .RN(n20700), .Q(n5293), 
        .QN(n19206) );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(n4301), .CK(CLK), .RN(n20745), .Q(n5292), 
        .QN(n19205) );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(n4300), .CK(CLK), .RN(n20701), .Q(n5291), 
        .QN(n19204) );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(n4299), .CK(CLK), .RN(n20724), .Q(n5290), 
        .QN(n19203) );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(n4298), .CK(CLK), .RN(n20728), .Q(n19578), .QN(n8685) );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(n4297), .CK(CLK), .RN(n20715), .Q(n19586), .QN(n8688) );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(n4296), .CK(CLK), .RN(n20698), .Q(n19577), .QN(n8687) );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(n4295), .CK(CLK), .RN(n20706), .Q(n19576), .QN(n8684) );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(n4294), .CK(CLK), .RN(n20712), .Q(n19585), .QN(n8683) );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(n4293), .CK(CLK), .RN(n20692), .Q(n19575), .QN(n8686) );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(n4292), .CK(CLK), .RN(n20708), .Q(n19574), .QN(n8682) );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(n4291), .CK(CLK), .RN(n20699), .Q(n19573), .QN(n8681) );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(n4290), .CK(CLK), .RN(n20741), .Q(n19584), .QN(n8680) );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(n4289), .CK(CLK), .RN(n20700), .Q(n19572), .QN(n8679) );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(n4288), .CK(CLK), .RN(n20722), .Q(n19571), .QN(n8678) );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(n4287), .CK(CLK), .RN(n20719), .Q(n19570), .QN(n8677) );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(n4286), .CK(CLK), .RN(n20727), .Q(n19569), .QN(n8670) );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(n4285), .CK(CLK), .RN(n20742), .Q(n19568), .QN(n8669) );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(n4284), .CK(CLK), .RN(n20704), .Q(n19567), .QN(n8676) );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(n4283), .CK(CLK), .RN(n20735), .Q(n19583), .QN(n8668) );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(n4282), .CK(CLK), .RN(n20738), .Q(n19566), .QN(n8667) );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(n4281), .CK(CLK), .RN(n20701), .Q(n19565), .QN(n8675) );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(n4280), .CK(CLK), .RN(n20701), .Q(n19564), .QN(n8674) );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(n4279), .CK(CLK), .RN(n20702), .Q(n19582), .QN(n8673) );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(n4278), .CK(CLK), .RN(n20697), .Q(n19563), .QN(n8672) );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(n4277), .CK(CLK), .RN(n20716), .Q(n19562), .QN(n8666) );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(n4276), .CK(CLK), .RN(n20717), .Q(n19581), 
        .QN(n8665) );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(n4275), .CK(CLK), .RN(n20733), .Q(n19561), 
        .QN(n8671) );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(n4274), .CK(CLK), .RN(n20745), .Q(n19560), 
        .QN(n8664) );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(n4273), .CK(CLK), .RN(n20697), .Q(n19559), 
        .QN(n8663) );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(n4272), .CK(CLK), .RN(n20713), .Q(n19580), 
        .QN(n8662) );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(n4271), .CK(CLK), .RN(n20696), .Q(n19558), 
        .QN(n8661) );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(n4270), .CK(CLK), .RN(n20743), .Q(n19557), 
        .QN(n8660) );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(n4269), .CK(CLK), .RN(n20728), .Q(n19556), 
        .QN(n8659) );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(n4268), .CK(CLK), .RN(n20707), .Q(n19579), 
        .QN(n8658) );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(n4267), .CK(CLK), .RN(n20709), .Q(n19555), 
        .QN(n8657) );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(n4266), .CK(CLK), .RN(n20728), .Q(n17608), .QN(n8485) );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(n4265), .CK(CLK), .RN(n20718), .Q(n17616), .QN(n8484) );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(n4264), .CK(CLK), .RN(n20714), .Q(n17607), .QN(n8483) );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(n4263), .CK(CLK), .RN(n20740), .Q(n17606), .QN(n8481) );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(n4262), .CK(CLK), .RN(n20728), .Q(n17615), .QN(n8480) );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(n4261), .CK(CLK), .RN(n20722), .Q(n17605), .QN(n8482) );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(n4260), .CK(CLK), .RN(n20726), .Q(n17604), .QN(n8479) );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(n4259), .CK(CLK), .RN(n20699), .Q(n17603), .QN(n8478) );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(n4258), .CK(CLK), .RN(n20741), .Q(n17614), .QN(n8477) );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(n4257), .CK(CLK), .RN(n20714), .Q(n17602), .QN(n8476) );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(n4256), .CK(CLK), .RN(n20699), .Q(n17601), .QN(n8475) );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(n4255), .CK(CLK), .RN(n20724), .Q(n17600), .QN(n8474) );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(n4254), .CK(CLK), .RN(n20741), .Q(n17599), .QN(n8458) );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(n4253), .CK(CLK), .RN(n20701), .Q(n17598), .QN(n8472) );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(n4252), .CK(CLK), .RN(n20737), .Q(n17597), .QN(n8473) );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(n4251), .CK(CLK), .RN(n20735), .Q(n17613), .QN(n8471) );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(n4250), .CK(CLK), .RN(n20738), .Q(n17596), .QN(n8470) );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(n4249), .CK(CLK), .RN(n20736), .Q(n17595), .QN(n8469) );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(n4248), .CK(CLK), .RN(n20701), .Q(n17594), .QN(n8466) );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(n4247), .CK(CLK), .RN(n20728), .Q(n17612), .QN(n8465) );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(n4246), .CK(CLK), .RN(n20720), .Q(n17593), .QN(n8468) );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(n4245), .CK(CLK), .RN(n20709), .Q(n17592), .QN(n8464) );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(n4244), .CK(CLK), .RN(n20740), .Q(n17611), 
        .QN(n8463) );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(n4243), .CK(CLK), .RN(n20733), .Q(n17591), 
        .QN(n8467) );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(n4242), .CK(CLK), .RN(n20745), .Q(n17590), 
        .QN(n8462) );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(n4241), .CK(CLK), .RN(n20697), .Q(n17589), 
        .QN(n8461) );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(n4240), .CK(CLK), .RN(n20712), .Q(n17610), 
        .QN(n8460) );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(n4239), .CK(CLK), .RN(n20696), .Q(n17588), 
        .QN(n8457) );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(n4238), .CK(CLK), .RN(n20691), .Q(n17587), 
        .QN(n8456) );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(n4237), .CK(CLK), .RN(n20703), .Q(n17586), 
        .QN(n8459) );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(n4236), .CK(CLK), .RN(n20694), .Q(n17609), 
        .QN(n8455) );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(n4235), .CK(CLK), .RN(n20720), .Q(n17585), 
        .QN(n8454) );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(n4234), .CK(CLK), .RN(n20728), .Q(n5289), 
        .QN(n19650) );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(n4233), .CK(CLK), .RN(n20715), .Q(n5288), 
        .QN(n19649) );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(n4232), .CK(CLK), .RN(n20714), .Q(n5287), 
        .QN(n19648) );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(n4231), .CK(CLK), .RN(n20706), .Q(n5286), 
        .QN(n19647) );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(n4230), .CK(CLK), .RN(n20728), .Q(n5628), 
        .QN(n19646) );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(n4229), .CK(CLK), .RN(n20722), .Q(n5627), 
        .QN(n19645) );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(n4228), .CK(CLK), .RN(n20726), .Q(n5626), 
        .QN(n19644) );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(n4227), .CK(CLK), .RN(n20699), .Q(n5625), 
        .QN(n19643) );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(n4226), .CK(CLK), .RN(n20734), .Q(n5624), 
        .QN(n19642) );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(n4225), .CK(CLK), .RN(n20714), .Q(n5623), 
        .QN(n19641) );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(n4224), .CK(CLK), .RN(n20737), .Q(n5622), 
        .QN(n19640) );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(n4223), .CK(CLK), .RN(n20711), .Q(n5621), 
        .QN(n19639) );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(n4222), .CK(CLK), .RN(n20727), .Q(n5285), 
        .QN(n19638) );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(n4221), .CK(CLK), .RN(n20704), .Q(n5284), 
        .QN(n19637) );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(n4220), .CK(CLK), .RN(n20737), .Q(n5283), 
        .QN(n19636) );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(n4219), .CK(CLK), .RN(n20730), .Q(n5282), 
        .QN(n19635) );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(n4218), .CK(CLK), .RN(n20727), .Q(n5281), 
        .QN(n19634) );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(n4217), .CK(CLK), .RN(n20722), .Q(n5280), 
        .QN(n19633) );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(n4216), .CK(CLK), .RN(n20701), .Q(n5279), 
        .QN(n19632) );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(n4215), .CK(CLK), .RN(n20702), .Q(n5278), 
        .QN(n19631) );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(n4214), .CK(CLK), .RN(n20744), .Q(n5277), 
        .QN(n19630) );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(n4213), .CK(CLK), .RN(n20709), .Q(n5276), 
        .QN(n19629) );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(n4212), .CK(CLK), .RN(n20740), .Q(n5275), 
        .QN(n19628) );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(n4211), .CK(CLK), .RN(n20733), .Q(n5274), 
        .QN(n19627) );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(n4210), .CK(CLK), .RN(n20745), .Q(n5273), 
        .QN(n19626) );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(n4209), .CK(CLK), .RN(n20697), .Q(n5272), 
        .QN(n19625) );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(n4208), .CK(CLK), .RN(n20712), .Q(n5271), 
        .QN(n19624) );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(n4207), .CK(CLK), .RN(n20707), .Q(n5270), 
        .QN(n19623) );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(n4206), .CK(CLK), .RN(n20716), .Q(n5000), 
        .QN(n19622) );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(n4205), .CK(CLK), .RN(n20733), .Q(n4999), 
        .QN(n19621) );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(n4204), .CK(CLK), .RN(n20736), .Q(n4998), 
        .QN(n19620) );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(n4203), .CK(CLK), .RN(n20709), .Q(n4997), 
        .QN(n19619) );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(n4202), .CK(CLK), .RN(n20728), .Q(n5070), 
        .QN(n19378) );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(n4201), .CK(CLK), .RN(n20718), .Q(n5069), 
        .QN(n19384) );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(n4200), .CK(CLK), .RN(n20714), .Q(n5068), 
        .QN(n19392) );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(n4199), .CK(CLK), .RN(n20740), .Q(n5067), 
        .QN(n19377) );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(n4198), .CK(CLK), .RN(n20732), .Q(n5336), 
        .QN(n19383) );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(n4197), .CK(CLK), .RN(n20729), .Q(n5334), 
        .QN(n19391) );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(n4196), .CK(CLK), .RN(n20707), .Q(n5204), 
        .QN(n19376) );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(n4195), .CK(CLK), .RN(n20698), .Q(n5202), 
        .QN(n19375) );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(n4194), .CK(CLK), .RN(n20741), .Q(n5200), 
        .QN(n19394) );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(n4193), .CK(CLK), .RN(n20714), .Q(n5198), 
        .QN(n19374) );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(n4192), .CK(CLK), .RN(n20692), .Q(n5473), 
        .QN(n19373) );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(n4191), .CK(CLK), .RN(n20710), .Q(n5472), 
        .QN(n19390) );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(n4190), .CK(CLK), .RN(n20727), .Q(n5066), 
        .QN(n19372) );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(n4189), .CK(CLK), .RN(n20743), .Q(n5065), 
        .QN(n19371) );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(n4188), .CK(CLK), .RN(n20720), .Q(n5064), 
        .QN(n19389) );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(n4187), .CK(CLK), .RN(n20694), .Q(n5063), 
        .QN(n19382) );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(n4186), .CK(CLK), .RN(n20729), .Q(n5062), 
        .QN(n19370) );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(n4185), .CK(CLK), .RN(n20715), .Q(n5061), 
        .QN(n19388) );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(n4184), .CK(CLK), .RN(n20743), .Q(n5060), 
        .QN(n19369) );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(n4183), .CK(CLK), .RN(n20694), .Q(n5059), 
        .QN(n19381) );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(n4182), .CK(CLK), .RN(n20697), .Q(n5058), 
        .QN(n19387) );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(n4181), .CK(CLK), .RN(n20709), .Q(n5057), 
        .QN(n19368) );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(n4180), .CK(CLK), .RN(n20716), .Q(n5056), 
        .QN(n19380) );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(n4179), .CK(CLK), .RN(n20733), .Q(n5055), 
        .QN(n19386) );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(n4178), .CK(CLK), .RN(n20742), .Q(n5054), 
        .QN(n19367) );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(n4177), .CK(CLK), .RN(n20697), .Q(n5053), 
        .QN(n19366) );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(n4176), .CK(CLK), .RN(n20712), .Q(n5052), 
        .QN(n19393) );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(n4175), .CK(CLK), .RN(n20707), .Q(n5051), 
        .QN(n19365) );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(n4174), .CK(CLK), .RN(n20720), .Q(n5050), 
        .QN(n19364) );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(n4173), .CK(CLK), .RN(n20717), .Q(n5049), 
        .QN(n19385) );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(n4172), .CK(CLK), .RN(n20721), .Q(n5048), 
        .QN(n19379) );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(n4171), .CK(CLK), .RN(n20724), .Q(n5047), 
        .QN(n19363) );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(n4170), .CK(CLK), .RN(n20739), .Q(n5215), 
        .QN(n19090) );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(n4169), .CK(CLK), .RN(n20724), .Q(n5214), 
        .QN(n19096) );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(n4168), .CK(CLK), .RN(n20697), .Q(n5213), 
        .QN(n19104) );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(n4167), .CK(CLK), .RN(n20742), .Q(n5212), 
        .QN(n19089) );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(n4166), .CK(CLK), .RN(n20704), .Q(n5211), 
        .QN(n19095) );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(n4165), .CK(CLK), .RN(n20709), .Q(n5210), 
        .QN(n19103) );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(n4164), .CK(CLK), .RN(n20708), .Q(n5209), 
        .QN(n19088) );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(n4163), .CK(CLK), .RN(n20726), .Q(n5208), 
        .QN(n19087) );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(n4162), .CK(CLK), .RN(n20734), .Q(n5207), 
        .QN(n19106) );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(n4161), .CK(CLK), .RN(n20719), .Q(n5206), 
        .QN(n19086) );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(n4160), .CK(CLK), .RN(n20692), .Q(n5265), 
        .QN(n19085) );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(n4159), .CK(CLK), .RN(n20710), .Q(n5264), 
        .QN(n19102) );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(n4158), .CK(CLK), .RN(n20727), .Q(n5263), 
        .QN(n19084) );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(n4157), .CK(CLK), .RN(n20737), .Q(n5262), 
        .QN(n19083) );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(n4156), .CK(CLK), .RN(n20724), .Q(n5261), 
        .QN(n19101) );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(n4155), .CK(CLK), .RN(n20702), .Q(n5260), 
        .QN(n19094) );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(n4154), .CK(CLK), .RN(n20730), .Q(n5259), 
        .QN(n19082) );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(n4153), .CK(CLK), .RN(n20712), .Q(n5258), 
        .QN(n19100) );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(n4152), .CK(CLK), .RN(n20743), .Q(n5257), 
        .QN(n19081) );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(n4151), .CK(CLK), .RN(n20694), .Q(n5256), 
        .QN(n19093) );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(n4150), .CK(CLK), .RN(n20743), .Q(n5255), 
        .QN(n19099) );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(n4149), .CK(CLK), .RN(n20706), .Q(n5254), 
        .QN(n19080) );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(n4148), .CK(CLK), .RN(n20710), .Q(n5253), 
        .QN(n19092) );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(n4147), .CK(CLK), .RN(n20733), .Q(n5252), 
        .QN(n19098) );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(n4146), .CK(CLK), .RN(n20742), .Q(n5251), 
        .QN(n19079) );
  DFFR_X1 \REGISTERS_reg[8][6]  ( .D(n4145), .CK(CLK), .RN(n20718), .Q(n5250), 
        .QN(n19078) );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(n4144), .CK(CLK), .RN(n20718), .Q(n5249), 
        .QN(n19105) );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(n4143), .CK(CLK), .RN(n20734), .Q(n5248), 
        .QN(n19077) );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(n4142), .CK(CLK), .RN(n20739), .Q(n5247), 
        .QN(n19076) );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(n4141), .CK(CLK), .RN(n20725), .Q(n5246), 
        .QN(n19097) );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(n4140), .CK(CLK), .RN(n20742), .Q(n5245), 
        .QN(n19091) );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(n4139), .CK(CLK), .RN(n20738), .Q(n5244), 
        .QN(n19075) );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(n4138), .CK(CLK), .RN(n20728), .Q(n19522), .QN(n4895) );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(n4137), .CK(CLK), .RN(n20709), .Q(n19521), .QN(n4894) );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(n4136), .CK(CLK), .RN(n20704), .Q(n19520), .QN(n4893) );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(n4135), .CK(CLK), .RN(n20742), .Q(n19519), .QN(n4892) );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(n4134), .CK(CLK), .RN(n20712), .Q(n19518), .QN(n4891) );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(n4133), .CK(CLK), .RN(n20722), .Q(n19517), .QN(n4890) );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(n4132), .CK(CLK), .RN(n20708), .Q(n19516), .QN(n4889) );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(n4131), .CK(CLK), .RN(n20698), .Q(n19515), .QN(n5150) );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(n4130), .CK(CLK), .RN(n20718), .Q(n19514), .QN(n5149) );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(n4129), .CK(CLK), .RN(n20725), .Q(n19513), .QN(n5148) );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(n4128), .CK(CLK), .RN(n20693), .Q(n19512), .QN(n5147) );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(n4127), .CK(CLK), .RN(n20724), .Q(n19511), .QN(n5146) );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(n4126), .CK(CLK), .RN(n20698), .Q(n19510), .QN(n5145) );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(n4125), .CK(CLK), .RN(n20731), .Q(n19509), .QN(n5144) );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(n4124), .CK(CLK), .RN(n20716), .Q(n19508), .QN(n5143) );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(n4123), .CK(CLK), .RN(n20702), .Q(n19507), .QN(n5142) );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(n4122), .CK(CLK), .RN(n20719), .Q(n19506), .QN(n5141) );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(n4121), .CK(CLK), .RN(n20712), .Q(n19505), .QN(n5140) );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(n4120), .CK(CLK), .RN(n20730), .Q(n19504), .QN(n5139) );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(n4119), .CK(CLK), .RN(n20743), .Q(n19503), .QN(n5138) );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(n4118), .CK(CLK), .RN(n20723), .Q(n19502), .QN(n5137) );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(n4117), .CK(CLK), .RN(n20715), .Q(n19501), .QN(n5136) );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(n4116), .CK(CLK), .RN(n20718), .Q(n19500), 
        .QN(n5135) );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(n4115), .CK(CLK), .RN(n20735), .Q(n19499), 
        .QN(n5134) );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(n4114), .CK(CLK), .RN(n20742), .Q(n19498), 
        .QN(n5133) );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(n4113), .CK(CLK), .RN(n20718), .Q(n19497), 
        .QN(n5132) );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(n4112), .CK(CLK), .RN(n20725), .Q(n19496), 
        .QN(n5131) );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(n4111), .CK(CLK), .RN(n20717), .Q(n19495), 
        .QN(n5130) );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(n4110), .CK(CLK), .RN(n20739), .Q(n19494), 
        .QN(n5129) );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(n4109), .CK(CLK), .RN(n20729), .Q(n19493), 
        .QN(n5128) );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(n4108), .CK(CLK), .RN(n20725), .Q(n19492), 
        .QN(n5127) );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(n4107), .CK(CLK), .RN(n20737), .Q(n19491), 
        .QN(n5126) );
  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(n4106), .CK(CLK), .RN(n20726), .Q(n5232), .QN(n18978) );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(n4105), .CK(CLK), .RN(n20726), .Q(n5231), .QN(n18977) );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(n4104), .CK(CLK), .RN(n20740), .Q(n5221), .QN(n18976) );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(n4103), .CK(CLK), .RN(n20744), .Q(n5230), .QN(n18975) );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(n4102), .CK(CLK), .RN(n20707), .Q(n5229), .QN(n18974) );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(n4101), .CK(CLK), .RN(n20703), .Q(n5220), .QN(n18973) );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(n4100), .CK(CLK), .RN(n20720), .Q(n5228), .QN(n18972) );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(n4099), .CK(CLK), .RN(n20710), .Q(n5227), .QN(n18971) );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(n4098), .CK(CLK), .RN(n20734), .Q(n5219), .QN(n18970) );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(n4097), .CK(CLK), .RN(n20701), .Q(n5226), .QN(n18969) );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(n4096), .CK(CLK), .RN(n20738), .Q(n5269), .QN(n18968) );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(n4095), .CK(CLK), .RN(n20719), .Q(n5268), .QN(n18967) );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(n4094), .CK(CLK), .RN(n20715), .Q(n5267), .QN(n18966) );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(n4093), .CK(CLK), .RN(n20696), .Q(n5266), .QN(n18965) );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(n4092), .CK(CLK), .RN(n20691), .Q(n5218), .QN(n18964) );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(n4091), .CK(CLK), .RN(n20746), .Q(n5225), .QN(n18963) );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(n4090), .CK(CLK), .RN(n20703), .Q(n5224), .QN(n18962) );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(n4089), .CK(CLK), .RN(n20735), .Q(n5217), .QN(n18961) );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(n4088), .CK(CLK), .RN(n20699), .Q(n5223), .QN(n18960) );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(n4087), .CK(CLK), .RN(n20710), .Q(n5222), .QN(n18959) );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(n4086), .CK(CLK), .RN(n20710), .Q(n5216), .QN(n18958) );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(n4085), .CK(CLK), .RN(n20692), .Q(n5243), .QN(n18957) );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(n4084), .CK(CLK), .RN(n20710), .Q(n5242), 
        .QN(n18956) );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(n4083), .CK(CLK), .RN(n20719), .Q(n5241), 
        .QN(n18955) );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(n4082), .CK(CLK), .RN(n20725), .Q(n5240), 
        .QN(n18954) );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(n4081), .CK(CLK), .RN(n20708), .Q(n5239), 
        .QN(n18953) );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(n4080), .CK(CLK), .RN(n20712), .Q(n5238), 
        .QN(n18952) );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(n4079), .CK(CLK), .RN(n20706), .Q(n5237), 
        .QN(n18951) );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(n4078), .CK(CLK), .RN(n20733), .Q(n5236), 
        .QN(n18950) );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(n4077), .CK(CLK), .RN(n20739), .Q(n5235), 
        .QN(n18949) );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(n4076), .CK(CLK), .RN(n20733), .Q(n5234), 
        .QN(n18948) );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(n4075), .CK(CLK), .RN(n20692), .Q(n5233), 
        .QN(n18947) );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(n4074), .CK(CLK), .RN(n20704), .Q(n4834), .QN(n19778) );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(n4073), .CK(CLK), .RN(n20732), .Q(n4833), .QN(n19777) );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(n4072), .CK(CLK), .RN(n20722), .Q(n4832), .QN(n19776) );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(n4071), .CK(CLK), .RN(n20744), .Q(n4831), .QN(n19775) );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(n4070), .CK(CLK), .RN(n20735), .Q(n4830), .QN(n19774) );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(n4069), .CK(CLK), .RN(n20737), .Q(n4829), .QN(n19773) );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(n4068), .CK(CLK), .RN(n20692), .Q(n4828), .QN(n19772) );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(n4067), .CK(CLK), .RN(n20737), .Q(n4827), .QN(n19771) );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(n4066), .CK(CLK), .RN(n20734), .Q(n4826), .QN(n19770) );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(n4065), .CK(CLK), .RN(n20734), .Q(n4825), .QN(n19769) );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(n4064), .CK(CLK), .RN(n20703), .Q(n4824), .QN(n19768) );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(n4063), .CK(CLK), .RN(n20719), .Q(n4823), .QN(n19767) );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(n4062), .CK(CLK), .RN(n20715), .Q(n4822), .QN(n19766) );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(n4061), .CK(CLK), .RN(n20696), .Q(n4821), .QN(n19765) );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(n4060), .CK(CLK), .RN(n20703), .Q(n4820), .QN(n19764) );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(n4059), .CK(CLK), .RN(n20702), .Q(n4819), .QN(n19763) );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(n4058), .CK(CLK), .RN(n20728), .Q(n4818), .QN(n19762) );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(n4057), .CK(CLK), .RN(n20746), .Q(n4817), .QN(n19761) );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(n4056), .CK(CLK), .RN(n20693), .Q(n4816), .QN(n19760) );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(n4055), .CK(CLK), .RN(n20716), .Q(n4815), .QN(n19759) );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(n4054), .CK(CLK), .RN(n20727), .Q(n4814), .QN(n19758) );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(n4053), .CK(CLK), .RN(n20692), .Q(n4813), .QN(n19757) );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(n4052), .CK(CLK), .RN(n20745), .Q(n4812), 
        .QN(n19756) );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(n4051), .CK(CLK), .RN(n20702), .Q(n4811), 
        .QN(n19755) );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(n4050), .CK(CLK), .RN(n20725), .Q(n4810), 
        .QN(n19754) );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(n4049), .CK(CLK), .RN(n20733), .Q(n4809), 
        .QN(n19753) );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(n4048), .CK(CLK), .RN(n20712), .Q(n4808), 
        .QN(n19752) );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(n4047), .CK(CLK), .RN(n20706), .Q(n4807), 
        .QN(n19751) );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(n4046), .CK(CLK), .RN(n20743), .Q(n4806), 
        .QN(n19750) );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(n4045), .CK(CLK), .RN(n20712), .Q(n4805), 
        .QN(n19749) );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(n4044), .CK(CLK), .RN(n20733), .Q(n4804), 
        .QN(n19748) );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(n4043), .CK(CLK), .RN(n20737), .Q(n4803), 
        .QN(n19747) );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(n4042), .CK(CLK), .RN(n20742), .Q(
        n19010), .QN(n5602) );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(n4041), .CK(CLK), .RN(n20709), .Q(
        n19009), .QN(n5601) );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(n4040), .CK(CLK), .RN(n20691), .Q(
        n19008), .QN(n5600) );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(n4039), .CK(CLK), .RN(n20742), .Q(
        n19007), .QN(n5599) );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(n4038), .CK(CLK), .RN(n20705), .Q(
        n19006), .QN(n5598) );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(n4037), .CK(CLK), .RN(n20722), .Q(
        n19005), .QN(n5597) );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(n4036), .CK(CLK), .RN(n20699), .Q(
        n19004), .QN(n5596) );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(n4035), .CK(CLK), .RN(n20698), .Q(
        n19003), .QN(n5595) );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(n4034), .CK(CLK), .RN(n20734), .Q(
        n19002), .QN(n5478) );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(n4033), .CK(CLK), .RN(n20700), .Q(
        n19001), .QN(n5594) );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(n4032), .CK(CLK), .RN(n20693), .Q(
        n19000), .QN(n5593) );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(n4031), .CK(CLK), .RN(n20724), .Q(
        n18999), .QN(n5592) );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(n4030), .CK(CLK), .RN(n20713), .Q(
        n18998), .QN(n5591) );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(n4029), .CK(CLK), .RN(n20693), .Q(
        n18997), .QN(n5590) );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(n4028), .CK(CLK), .RN(n20716), .Q(
        n18996), .QN(n5589) );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(n4027), .CK(CLK), .RN(n20706), .Q(
        n18995), .QN(n5588) );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(n4026), .CK(CLK), .RN(n20712), .Q(
        n18994), .QN(n5587) );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(n4025), .CK(CLK), .RN(n20736), .Q(
        n18993), .QN(n5586) );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(n4024), .CK(CLK), .RN(n20739), .Q(
        n18992), .QN(n5585) );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(n4023), .CK(CLK), .RN(n20721), .Q(
        n18991), .QN(n5584) );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(n4022), .CK(CLK), .RN(n20713), .Q(
        n18990), .QN(n5583) );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(n4021), .CK(CLK), .RN(n20741), .Q(
        n18989), .QN(n5582) );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(n4020), .CK(CLK), .RN(n20743), .Q(n18988), .QN(n5581) );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(n4019), .CK(CLK), .RN(n20706), .Q(n18987), .QN(n5580) );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(n4018), .CK(CLK), .RN(n20717), .Q(n18986), .QN(n5579) );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(n4017), .CK(CLK), .RN(n20711), .Q(n18985), .QN(n5578) );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(n4016), .CK(CLK), .RN(n20696), .Q(n18984), .QN(n5577) );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(n4015), .CK(CLK), .RN(n20717), .Q(n18983), .QN(n5576) );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(n4014), .CK(CLK), .RN(n20739), .Q(n18982), .QN(n5575) );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(n4013), .CK(CLK), .RN(n20729), .Q(n18981), .QN(n5574) );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(n4012), .CK(CLK), .RN(n20691), .Q(n18980), .QN(n5573) );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(n4011), .CK(CLK), .RN(n20724), .Q(n18979), .QN(n5572) );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(n4010), .CK(CLK), .RN(n20730), .Q(n5866), .QN(n19320) );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(n4009), .CK(CLK), .RN(n20709), .Q(n5865), .QN(n19319) );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(n4008), .CK(CLK), .RN(n20704), .Q(n5864), .QN(n19330) );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(n4007), .CK(CLK), .RN(n20721), .Q(n5863), .QN(n19318) );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(n4006), .CK(CLK), .RN(n20705), .Q(n5862), .QN(n19317) );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(n4005), .CK(CLK), .RN(n20722), .Q(n5861), .QN(n19329) );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(n4004), .CK(CLK), .RN(n20720), .Q(n5860), .QN(n19316) );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(n4003), .CK(CLK), .RN(n20698), .Q(n5859), .QN(n19315) );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(n4002), .CK(CLK), .RN(n20741), .Q(n5858), .QN(n19328) );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(n4001), .CK(CLK), .RN(n20725), .Q(n5857), .QN(n19314) );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(n4000), .CK(CLK), .RN(n20693), .Q(n5856), .QN(n19313) );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(n3999), .CK(CLK), .RN(n20729), .Q(n5855), .QN(n19327) );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(n3998), .CK(CLK), .RN(n20733), .Q(n5854), .QN(n19312) );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(n3997), .CK(CLK), .RN(n20694), .Q(n5853), .QN(n19311) );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(n3996), .CK(CLK), .RN(n20730), .Q(n5852), .QN(n19326) );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(n3995), .CK(CLK), .RN(n20706), .Q(n5851), .QN(n19310) );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(n3994), .CK(CLK), .RN(n20730), .Q(n5850), .QN(n19309) );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(n3993), .CK(CLK), .RN(n20712), .Q(n5849), .QN(n19325) );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(n3992), .CK(CLK), .RN(n20716), .Q(n5848), .QN(n19308) );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(n3991), .CK(CLK), .RN(n20720), .Q(n5847), .QN(n19307) );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(n3990), .CK(CLK), .RN(n20713), .Q(n5846), .QN(n19324) );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(n3989), .CK(CLK), .RN(n20710), .Q(n5845), .QN(n19306) );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(n3988), .CK(CLK), .RN(n20743), .Q(n5844), 
        .QN(n19305) );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(n3987), .CK(CLK), .RN(n20706), .Q(n5843), 
        .QN(n19323) );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(n3986), .CK(CLK), .RN(n20742), .Q(n5842), 
        .QN(n19304) );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(n3985), .CK(CLK), .RN(n20703), .Q(n5841), 
        .QN(n19303) );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(n3984), .CK(CLK), .RN(n20729), .Q(n5840), 
        .QN(n19322) );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(n3983), .CK(CLK), .RN(n20720), .Q(n5839), 
        .QN(n19302) );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(n3982), .CK(CLK), .RN(n20710), .Q(n5838), 
        .QN(n19301) );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(n3981), .CK(CLK), .RN(n20729), .Q(n5837), 
        .QN(n19321) );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(n3980), .CK(CLK), .RN(n20724), .Q(n5836), 
        .QN(n19300) );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(n3979), .CK(CLK), .RN(n20732), .Q(n5835), 
        .QN(n19299) );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(n3978), .CK(CLK), .RN(n20716), .Q(n5036), .QN(n19442) );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(n3977), .CK(CLK), .RN(n20737), .Q(n5035), .QN(n19448) );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(n3976), .CK(CLK), .RN(n20691), .Q(n5046), .QN(n19456) );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(n3975), .CK(CLK), .RN(n20721), .Q(n5034), .QN(n19441) );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(n3974), .CK(CLK), .RN(n20728), .Q(n5033), .QN(n19447) );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(n3973), .CK(CLK), .RN(n20737), .Q(n5045), .QN(n19455) );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(n3972), .CK(CLK), .RN(n20720), .Q(n5032), .QN(n19440) );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(n3971), .CK(CLK), .RN(n20737), .Q(n5031), .QN(n19439) );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(n3970), .CK(CLK), .RN(n20741), .Q(n5044), .QN(n19458) );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(n3969), .CK(CLK), .RN(n20714), .Q(n5030), .QN(n19438) );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(n3968), .CK(CLK), .RN(n20737), .Q(n5029), .QN(n19437) );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(n3967), .CK(CLK), .RN(n20705), .Q(n5043), .QN(n19454) );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(n3966), .CK(CLK), .RN(n20733), .Q(n5028), .QN(n19436) );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(n3965), .CK(CLK), .RN(n20743), .Q(n5027), .QN(n19435) );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(n3964), .CK(CLK), .RN(n20730), .Q(n5042), .QN(n19453) );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(n3963), .CK(CLK), .RN(n20713), .Q(n5026), .QN(n19446) );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(n3962), .CK(CLK), .RN(n20732), .Q(n5025), .QN(n19434) );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(n3961), .CK(CLK), .RN(n20694), .Q(n5041), .QN(n19452) );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(n3960), .CK(CLK), .RN(n20704), .Q(n5024), .QN(n19433) );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(n3959), .CK(CLK), .RN(n20695), .Q(n5023), .QN(n19445) );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(n3958), .CK(CLK), .RN(n20743), .Q(n5040), .QN(n19451) );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(n3957), .CK(CLK), .RN(n20741), .Q(n5022), .QN(n19432) );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(n3956), .CK(CLK), .RN(n20695), .Q(n5021), 
        .QN(n19444) );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(n3955), .CK(CLK), .RN(n20706), .Q(n5039), 
        .QN(n19450) );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(n3954), .CK(CLK), .RN(n20742), .Q(n5020), 
        .QN(n19431) );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(n3953), .CK(CLK), .RN(n20739), .Q(n5019), 
        .QN(n19430) );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(n3952), .CK(CLK), .RN(n20699), .Q(n5038), 
        .QN(n19457) );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(n3951), .CK(CLK), .RN(n20732), .Q(n5018), 
        .QN(n19429) );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(n3950), .CK(CLK), .RN(n20704), .Q(n5017), 
        .QN(n19428) );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(n3949), .CK(CLK), .RN(n20729), .Q(n5037), 
        .QN(n19449) );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(n3948), .CK(CLK), .RN(n20740), .Q(n5016), 
        .QN(n19443) );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(n3947), .CK(CLK), .RN(n20738), .Q(n5015), 
        .QN(n19427) );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(n3946), .CK(CLK), .RN(n20721), .Q(
        n19610), .QN(n5571) );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(n3945), .CK(CLK), .RN(n20709), .Q(
        n19618), .QN(n5570) );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(n3944), .CK(CLK), .RN(n20691), .Q(
        n19609), .QN(n5569) );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(n3943), .CK(CLK), .RN(n20717), .Q(
        n19608), .QN(n5568) );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(n3942), .CK(CLK), .RN(n20706), .Q(
        n19617), .QN(n5567) );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(n3941), .CK(CLK), .RN(n20737), .Q(
        n19607), .QN(n5566) );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(n3940), .CK(CLK), .RN(n20720), .Q(
        n19606), .QN(n5565) );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(n3939), .CK(CLK), .RN(n20723), .Q(
        n19605), .QN(n5564) );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(n3938), .CK(CLK), .RN(n20708), .Q(
        n19616), .QN(n5477) );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(n3937), .CK(CLK), .RN(n20700), .Q(
        n19604), .QN(n5563) );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(n3936), .CK(CLK), .RN(n20722), .Q(
        n19603), .QN(n5562) );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(n3935), .CK(CLK), .RN(n20697), .Q(
        n19602), .QN(n5561) );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(n3934), .CK(CLK), .RN(n20717), .Q(
        n19601), .QN(n5560) );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(n3933), .CK(CLK), .RN(n20736), .Q(
        n19600), .QN(n5559) );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(n3932), .CK(CLK), .RN(n20716), .Q(
        n19599), .QN(n5558) );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(n3931), .CK(CLK), .RN(n20713), .Q(
        n19615), .QN(n5557) );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(n3930), .CK(CLK), .RN(n20692), .Q(
        n19598), .QN(n5556) );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(n3929), .CK(CLK), .RN(n20736), .Q(
        n19597), .QN(n5555) );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(n3928), .CK(CLK), .RN(n20721), .Q(
        n19596), .QN(n5554) );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(n3927), .CK(CLK), .RN(n20699), .Q(
        n19614), .QN(n5553) );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(n3926), .CK(CLK), .RN(n20707), .Q(
        n19595), .QN(n5552) );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(n3925), .CK(CLK), .RN(n20741), .Q(
        n19594), .QN(n5551) );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(n3924), .CK(CLK), .RN(n20695), .Q(n19613), .QN(n5550) );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(n3923), .CK(CLK), .RN(n20734), .Q(n19593), .QN(n5549) );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(n3922), .CK(CLK), .RN(n20730), .Q(n19592), .QN(n5548) );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(n3921), .CK(CLK), .RN(n20697), .Q(n19591), .QN(n5547) );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(n3920), .CK(CLK), .RN(n20713), .Q(n19612), .QN(n5546) );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(n3919), .CK(CLK), .RN(n20715), .Q(n19590), .QN(n5545) );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(n3918), .CK(CLK), .RN(n20734), .Q(n19589), .QN(n5544) );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(n3917), .CK(CLK), .RN(n20694), .Q(n19588), .QN(n5543) );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(n3916), .CK(CLK), .RN(n20724), .Q(n19611), .QN(n5542) );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(n3915), .CK(CLK), .RN(n20732), .Q(n19587), .QN(n5541) );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(n3914), .CK(CLK), .RN(n20736), .Q(
        n19546), .QN(n4888) );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(n3913), .CK(CLK), .RN(n20737), .Q(
        n19554), .QN(n4887) );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(n3912), .CK(CLK), .RN(n20707), .Q(
        n19545), .QN(n4886) );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(n3911), .CK(CLK), .RN(n20745), .Q(
        n19544), .QN(n4885) );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(n3910), .CK(CLK), .RN(n20710), .Q(
        n19553), .QN(n4884) );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(n3909), .CK(CLK), .RN(n20707), .Q(
        n19543), .QN(n4883) );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(n3908), .CK(CLK), .RN(n20709), .Q(
        n19542), .QN(n4882) );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(n3907), .CK(CLK), .RN(n20723), .Q(
        n19541), .QN(n4977) );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(n3906), .CK(CLK), .RN(n20741), .Q(
        n19552), .QN(n4975) );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(n3905), .CK(CLK), .RN(n20725), .Q(
        n19540), .QN(n4974) );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(n3904), .CK(CLK), .RN(n20696), .Q(
        n19539), .QN(n4973) );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(n3903), .CK(CLK), .RN(n20729), .Q(
        n19538), .QN(n4972) );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(n3902), .CK(CLK), .RN(n20733), .Q(
        n19537), .QN(n4971) );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(n3901), .CK(CLK), .RN(n20722), .Q(
        n19536), .QN(n4970) );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(n3900), .CK(CLK), .RN(n20730), .Q(
        n19535), .QN(n4969) );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(n3899), .CK(CLK), .RN(n20735), .Q(
        n19551), .QN(n4968) );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(n3898), .CK(CLK), .RN(n20721), .Q(
        n19534), .QN(n4967) );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(n3897), .CK(CLK), .RN(n20742), .Q(
        n19533), .QN(n4966) );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(n3896), .CK(CLK), .RN(n20722), .Q(
        n19532), .QN(n4965) );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(n3895), .CK(CLK), .RN(n20694), .Q(
        n19550), .QN(n4964) );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(n3894), .CK(CLK), .RN(n20718), .Q(
        n19531), .QN(n4963) );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(n3893), .CK(CLK), .RN(n20710), .Q(
        n19530), .QN(n4962) );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(n3892), .CK(CLK), .RN(n20695), .Q(n19549), .QN(n4961) );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(n3891), .CK(CLK), .RN(n20706), .Q(n19529), .QN(n4960) );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(n3890), .CK(CLK), .RN(n20734), .Q(n19528), .QN(n4959) );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(n3889), .CK(CLK), .RN(n20697), .Q(n19527), .QN(n4958) );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(n3888), .CK(CLK), .RN(n20691), .Q(n19548), .QN(n4957) );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(n3887), .CK(CLK), .RN(n20704), .Q(n19526), .QN(n4956) );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(n3886), .CK(CLK), .RN(n20709), .Q(n19525), .QN(n4955) );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(n3885), .CK(CLK), .RN(n20709), .Q(n19524), .QN(n4954) );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(n3884), .CK(CLK), .RN(n20736), .Q(n19547), .QN(n4953) );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(n3883), .CK(CLK), .RN(n20732), .Q(n19523), .QN(n4952) );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(n3882), .CK(CLK), .RN(n20736), .Q(
        n19170), .QN(n5540) );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(n3881), .CK(CLK), .RN(n20737), .Q(
        n19169), .QN(n5539) );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(n3880), .CK(CLK), .RN(n20729), .Q(
        n19168), .QN(n5538) );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(n3879), .CK(CLK), .RN(n20745), .Q(
        n19167), .QN(n5537) );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(n3878), .CK(CLK), .RN(n20744), .Q(
        n19166), .QN(n5536) );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(n3877), .CK(CLK), .RN(n20693), .Q(
        n19165), .QN(n5535) );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(n3876), .CK(CLK), .RN(n20709), .Q(
        n19164), .QN(n5534) );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(n3875), .CK(CLK), .RN(n20723), .Q(
        n19163), .QN(n5533) );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(n3874), .CK(CLK), .RN(n20725), .Q(
        n19162), .QN(n5476) );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(n3873), .CK(CLK), .RN(n20698), .Q(
        n19161), .QN(n5532) );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(n3872), .CK(CLK), .RN(n20696), .Q(
        n19160), .QN(n5531) );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(n3871), .CK(CLK), .RN(n20729), .Q(
        n19159), .QN(n5530) );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(n3870), .CK(CLK), .RN(n20718), .Q(
        n19158), .QN(n5529) );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(n3869), .CK(CLK), .RN(n20743), .Q(
        n19157), .QN(n5528) );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(n3868), .CK(CLK), .RN(n20716), .Q(
        n19156), .QN(n5527) );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(n3867), .CK(CLK), .RN(n20735), .Q(
        n19155), .QN(n5526) );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(n3866), .CK(CLK), .RN(n20714), .Q(
        n19154), .QN(n5525) );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(n3865), .CK(CLK), .RN(n20725), .Q(
        n19153), .QN(n5524) );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(n3864), .CK(CLK), .RN(n20721), .Q(
        n19152), .QN(n5523) );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(n3863), .CK(CLK), .RN(n20695), .Q(
        n19151), .QN(n5522) );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(n3862), .CK(CLK), .RN(n20731), .Q(
        n19150), .QN(n5521) );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(n3861), .CK(CLK), .RN(n20695), .Q(
        n19149), .QN(n5520) );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(n3860), .CK(CLK), .RN(n20695), .Q(n19148), .QN(n5519) );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(n3859), .CK(CLK), .RN(n20738), .Q(n19147), .QN(n5518) );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(n3858), .CK(CLK), .RN(n20740), .Q(n19146), .QN(n5517) );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(n3857), .CK(CLK), .RN(n20693), .Q(n19145), .QN(n5516) );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(n3856), .CK(CLK), .RN(n20691), .Q(n19144), .QN(n5515) );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(n3855), .CK(CLK), .RN(n20715), .Q(n19143), .QN(n5514) );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(n3854), .CK(CLK), .RN(n20704), .Q(n19142), .QN(n5513) );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(n3853), .CK(CLK), .RN(n20722), .Q(n19141), .QN(n5512) );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(n3852), .CK(CLK), .RN(n20736), .Q(n19140), .QN(n5511) );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(n3851), .CK(CLK), .RN(n20711), .Q(n19139), .QN(n5510) );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(n3850), .CK(CLK), .RN(n20736), .QN(
        n19138) );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(n3849), .CK(CLK), .RN(n20736), .QN(
        n19137) );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(n3848), .CK(CLK), .RN(n20707), .QN(
        n19136) );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(n3847), .CK(CLK), .RN(n20745), .QN(
        n19135) );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(n3846), .CK(CLK), .RN(n20744), .QN(
        n19134) );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(n3845), .CK(CLK), .RN(n20693), .QN(
        n19133) );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(n3844), .CK(CLK), .RN(n20731), .QN(
        n19132) );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(n3843), .CK(CLK), .RN(n20722), .QN(
        n19131) );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(n3842), .CK(CLK), .RN(n20737), .QN(
        n19130) );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(n3841), .CK(CLK), .RN(n20698), .QN(
        n19129) );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(n3840), .CK(CLK), .RN(n20696), .QN(
        n19128) );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(n3839), .CK(CLK), .RN(n20705), .QN(
        n19127) );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(n3838), .CK(CLK), .RN(n20697), .QN(
        n19126) );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(n3837), .CK(CLK), .RN(n20746), .QN(
        n19125) );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(n3836), .CK(CLK), .RN(n20700), .QN(
        n19124) );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(n3835), .CK(CLK), .RN(n20739), .QN(
        n19123) );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(n3834), .CK(CLK), .RN(n20740), .QN(
        n19122) );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(n3833), .CK(CLK), .RN(n20726), .QN(
        n19121) );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(n3832), .CK(CLK), .RN(n20738), .QN(
        n19120) );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(n3831), .CK(CLK), .RN(n20700), .QN(
        n19119) );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(n3830), .CK(CLK), .RN(n20735), .QN(
        n19118) );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(n3829), .CK(CLK), .RN(n20696), .QN(
        n19117) );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(n3828), .CK(CLK), .RN(n20695), .QN(
        n19116) );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(n3827), .CK(CLK), .RN(n20721), .QN(
        n19115) );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(n3826), .CK(CLK), .RN(n20706), .QN(
        n19114) );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(n3825), .CK(CLK), .RN(n20708), .QN(
        n19113) );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(n3824), .CK(CLK), .RN(n20725), .QN(
        n19112) );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(n3823), .CK(CLK), .RN(n20695), .QN(
        n19111) );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(n3822), .CK(CLK), .RN(n20704), .QN(
        n19110) );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(n3821), .CK(CLK), .RN(n20694), .QN(
        n19109) );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(n3820), .CK(CLK), .RN(n20701), .QN(
        n19108) );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(n3819), .CK(CLK), .RN(n20712), .QN(
        n19107) );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(n3818), .CK(CLK), .RN(n20719), .Q(n4802), .QN(n19258) );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(n3817), .CK(CLK), .RN(n20732), .Q(n4801), .QN(n19257) );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(n3816), .CK(CLK), .RN(n20714), .Q(n4800), .QN(n19256) );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(n3815), .CK(CLK), .RN(n20723), .Q(n4799), .QN(n19255) );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(n3814), .CK(CLK), .RN(n20740), .Q(n4842), .QN(n19266) );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(n3813), .CK(CLK), .RN(n20731), .Q(n4841), .QN(n19264) );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(n3812), .CK(CLK), .RN(n20720), .Q(n4840), .QN(n19263) );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(n3811), .CK(CLK), .RN(n20737), .Q(n4839), .QN(n19262) );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(n3810), .CK(CLK), .RN(n20704), .Q(n4838), .QN(n19265) );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(n3809), .CK(CLK), .RN(n20729), .Q(n4837), .QN(n19261) );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(n3808), .CK(CLK), .RN(n20703), .Q(n4836), .QN(n19260) );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(n3807), .CK(CLK), .RN(n20718), .Q(n4835), .QN(n19259) );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(n3806), .CK(CLK), .RN(n20715), .Q(n4798), .QN(n19254) );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(n3805), .CK(CLK), .RN(n20739), .Q(n4797), .QN(n19253) );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(n3804), .CK(CLK), .RN(n20730), .Q(n4796), .QN(n19252) );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(n3803), .CK(CLK), .RN(n20736), .Q(n4795), .QN(n19251) );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(n3802), .CK(CLK), .RN(n20728), .Q(n4794), .QN(n19250) );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(n3801), .CK(CLK), .RN(n20701), .Q(n4793), .QN(n19249) );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(n3800), .CK(CLK), .RN(n20706), .Q(n4792), .QN(n19248) );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(n3799), .CK(CLK), .RN(n20729), .Q(n4791), .QN(n19247) );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(n3798), .CK(CLK), .RN(n20727), .Q(n4790), .QN(n19246) );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(n3797), .CK(CLK), .RN(n20692), .Q(n4789), .QN(n19245) );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(n3796), .CK(CLK), .RN(n20699), .Q(n4788), 
        .QN(n19244) );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(n3795), .CK(CLK), .RN(n20740), .Q(n4787), 
        .QN(n19243) );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(n3794), .CK(CLK), .RN(n20713), .Q(n4786), 
        .QN(n19242) );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(n3793), .CK(CLK), .RN(n20693), .Q(n4785), 
        .QN(n19241) );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(n3792), .CK(CLK), .RN(n20726), .Q(n4784), 
        .QN(n19240) );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(n3791), .CK(CLK), .RN(n20706), .Q(n4783), 
        .QN(n19239) );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(n3790), .CK(CLK), .RN(n20701), .Q(n4782), 
        .QN(n19238) );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(n3789), .CK(CLK), .RN(n20745), .Q(n4781), 
        .QN(n19237) );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(n3788), .CK(CLK), .RN(n20713), .Q(n4780), 
        .QN(n19236) );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(n3787), .CK(CLK), .RN(n20711), .Q(n4779), 
        .QN(n19235) );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(n3786), .CK(CLK), .RN(n20736), .Q(
        n17488), .QN(n8517) );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(n3785), .CK(CLK), .RN(n20736), .Q(
        n17487), .QN(n8516) );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(n3784), .CK(CLK), .RN(n20707), .Q(
        n17486), .QN(n8515) );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(n3783), .CK(CLK), .RN(n20745), .Q(
        n17485), .QN(n8514) );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(n3782), .CK(CLK), .RN(n20744), .Q(
        n17484), .QN(n8513) );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(n3781), .CK(CLK), .RN(n20693), .Q(
        n17483), .QN(n8512) );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(n3780), .CK(CLK), .RN(n20732), .Q(
        n17482), .QN(n8511) );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(n3779), .CK(CLK), .RN(n20723), .Q(
        n17481), .QN(n8510) );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(n3778), .CK(CLK), .RN(n20731), .Q(
        n17480), .QN(n8509) );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(n3777), .CK(CLK), .RN(n20731), .Q(
        n17479), .QN(n8508) );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(n3776), .CK(CLK), .RN(n20703), .Q(
        n17478), .QN(n8507) );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(n3775), .CK(CLK), .RN(n20724), .Q(
        n17477), .QN(n8506) );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(n3774), .CK(CLK), .RN(n20715), .Q(
        n17476), .QN(n8505) );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(n3773), .CK(CLK), .RN(n20704), .Q(
        n17475), .QN(n8504) );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(n3772), .CK(CLK), .RN(n20736), .Q(
        n17474), .QN(n8503) );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(n3771), .CK(CLK), .RN(n20739), .Q(
        n17473), .QN(n8502) );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(n3770), .CK(CLK), .RN(n20738), .Q(
        n17472), .QN(n8501) );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(n3769), .CK(CLK), .RN(n20726), .Q(
        n17471), .QN(n8500) );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(n3768), .CK(CLK), .RN(n20701), .Q(
        n17470), .QN(n8499) );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(n3767), .CK(CLK), .RN(n20699), .Q(
        n17469), .QN(n8498) );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(n3766), .CK(CLK), .RN(n20739), .Q(
        n17468), .QN(n8497) );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(n3765), .CK(CLK), .RN(n20696), .Q(
        n17467), .QN(n8496) );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(n3764), .CK(CLK), .RN(n20745), .Q(n17466), .QN(n8495) );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(n3763), .CK(CLK), .RN(n20721), .Q(n17465), .QN(n8494) );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(n3762), .CK(CLK), .RN(n20740), .Q(n17464), .QN(n8493) );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(n3761), .CK(CLK), .RN(n20730), .Q(n17463), .QN(n8492) );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(n3760), .CK(CLK), .RN(n20725), .Q(n17462), .QN(n8491) );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(n3759), .CK(CLK), .RN(n20700), .Q(n17461), .QN(n8490) );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(n3758), .CK(CLK), .RN(n20738), .Q(n17460), .QN(n8489) );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(n3757), .CK(CLK), .RN(n20694), .Q(n17459), .QN(n8488) );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(n3756), .CK(CLK), .RN(n20730), .Q(n17458), .QN(n8487) );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(n3755), .CK(CLK), .RN(n20712), .Q(n17457), .QN(n8486) );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(n3754), .CK(CLK), .RN(n20694), .QN(
        n19074) );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(n3753), .CK(CLK), .RN(n20708), .QN(
        n19073) );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(n3752), .CK(CLK), .RN(n20729), .QN(
        n19072) );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(n3751), .CK(CLK), .RN(n20745), .QN(
        n19071) );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(n3750), .CK(CLK), .RN(n20744), .QN(
        n19070) );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(n3749), .CK(CLK), .RN(n20693), .QN(
        n19069) );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(n3748), .CK(CLK), .RN(n20731), .QN(
        n19068) );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(n3747), .CK(CLK), .RN(n20723), .QN(
        n19067) );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(n3746), .CK(CLK), .RN(n20731), .QN(
        n19066) );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(n3745), .CK(CLK), .RN(n20711), .QN(
        n19065) );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(n3744), .CK(CLK), .RN(n20717), .QN(
        n19064) );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(n3743), .CK(CLK), .RN(n20727), .QN(
        n19063) );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(n3742), .CK(CLK), .RN(n20733), .QN(
        n19062) );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(n3741), .CK(CLK), .RN(n20691), .QN(
        n19061) );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(n3740), .CK(CLK), .RN(n20699), .QN(
        n19060) );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(n3739), .CK(CLK), .RN(n20739), .QN(
        n19059) );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(n3738), .CK(CLK), .RN(n20714), .QN(
        n19058) );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(n3737), .CK(CLK), .RN(n20726), .QN(
        n19057) );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(n3736), .CK(CLK), .RN(n20709), .QN(
        n19056) );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(n3735), .CK(CLK), .RN(n20699), .QN(
        n19055) );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(n3734), .CK(CLK), .RN(n20707), .QN(
        n19054) );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(n3733), .CK(CLK), .RN(n20696), .QN(
        n19053) );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(n3732), .CK(CLK), .RN(n20707), .QN(
        n19052) );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(n3731), .CK(CLK), .RN(n20691), .QN(
        n19051) );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(n3730), .CK(CLK), .RN(n20740), .QN(
        n19050) );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(n3729), .CK(CLK), .RN(n20708), .QN(
        n19049) );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(n3728), .CK(CLK), .RN(n20725), .QN(
        n19048) );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(n3727), .CK(CLK), .RN(n20730), .QN(
        n19047) );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(n3726), .CK(CLK), .RN(n20738), .QN(
        n19046) );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(n3725), .CK(CLK), .RN(n20711), .QN(
        n19045) );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(n3724), .CK(CLK), .RN(n20707), .QN(
        n19044) );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(n3723), .CK(CLK), .RN(n20711), .QN(
        n19043) );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(n3722), .CK(CLK), .RN(n20719), .Q(n5175), .QN(n18906) );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(n3721), .CK(CLK), .RN(n20732), .Q(n5174), .QN(n18905) );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(n3720), .CK(CLK), .RN(n20698), .Q(n5173), .QN(n18904) );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(n3719), .CK(CLK), .RN(n20723), .Q(n5172), .QN(n18903) );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(n3718), .CK(CLK), .RN(n20740), .Q(n5455), .QN(n18914) );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(n3717), .CK(CLK), .RN(n20731), .Q(n5454), .QN(n18913) );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(n3716), .CK(CLK), .RN(n20701), .Q(n5453), .QN(n18912) );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(n3715), .CK(CLK), .RN(n20695), .Q(n5452), .QN(n18911) );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(n3714), .CK(CLK), .RN(n20705), .Q(n5451), .QN(n18910) );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(n3713), .CK(CLK), .RN(n20711), .Q(n5450), .QN(n18909) );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(n3712), .CK(CLK), .RN(n20717), .Q(n5449), .QN(n18908) );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(n3711), .CK(CLK), .RN(n20727), .Q(n5448), .QN(n18907) );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(n3710), .CK(CLK), .RN(n20716), .Q(n5171), .QN(n18902) );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(n3709), .CK(CLK), .RN(n20704), .Q(n5170), .QN(n18901) );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(n3708), .CK(CLK), .RN(n20703), .Q(n5169), .QN(n18900) );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(n3707), .CK(CLK), .RN(n20718), .Q(n5168), .QN(n18899) );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(n3706), .CK(CLK), .RN(n20733), .Q(n5167), .QN(n18898) );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(n3705), .CK(CLK), .RN(n20741), .Q(n5166), .QN(n18897) );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(n3704), .CK(CLK), .RN(n20743), .Q(n5165), .QN(n18896) );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(n3703), .CK(CLK), .RN(n20702), .Q(n5164), .QN(n18895) );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(n3702), .CK(CLK), .RN(n20727), .Q(n5163), .QN(n18894) );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(n3701), .CK(CLK), .RN(n20739), .Q(n5162), .QN(n18893) );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(n3700), .CK(CLK), .RN(n20715), .Q(n5161), 
        .QN(n18892) );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(n3699), .CK(CLK), .RN(n20719), .Q(n5160), 
        .QN(n18891) );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(n3698), .CK(CLK), .RN(n20711), .Q(n5159), 
        .QN(n18890) );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(n3697), .CK(CLK), .RN(n20740), .Q(n5158), 
        .QN(n18889) );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(n3696), .CK(CLK), .RN(n20735), .Q(n5157), 
        .QN(n18888) );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(n3695), .CK(CLK), .RN(n20725), .Q(n5156), 
        .QN(n18887) );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(n3694), .CK(CLK), .RN(n20700), .Q(n5155), 
        .QN(n18886) );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(n3693), .CK(CLK), .RN(n20745), .Q(n5154), 
        .QN(n18885) );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(n3692), .CK(CLK), .RN(n20713), .Q(n5153), 
        .QN(n18884) );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(n3691), .CK(CLK), .RN(n20712), .Q(n5152), 
        .QN(n18883) );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(n3690), .CK(CLK), .RN(n20695), .Q(n5736), .QN(n19298) );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(n3689), .CK(CLK), .RN(n20736), .Q(n5735), .QN(n19297) );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(n3688), .CK(CLK), .RN(n20705), .Q(n5734), .QN(n19296) );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(n3687), .CK(CLK), .RN(n20744), .Q(n5733), .QN(n19295) );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(n3686), .CK(CLK), .RN(n20744), .Q(n5744), .QN(n19294) );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(n3685), .CK(CLK), .RN(n20700), .Q(n5743), .QN(n19293) );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(n3684), .CK(CLK), .RN(n20702), .Q(n5742), .QN(n19292) );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(n3683), .CK(CLK), .RN(n20722), .Q(n5741), .QN(n19291) );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(n3682), .CK(CLK), .RN(n20731), .Q(n5740), .QN(n19290) );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(n3681), .CK(CLK), .RN(n20734), .Q(n5739), .QN(n19289) );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(n3680), .CK(CLK), .RN(n20717), .Q(n5738), .QN(n19288) );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(n3679), .CK(CLK), .RN(n20724), .Q(n5737), .QN(n19287) );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(n3678), .CK(CLK), .RN(n20744), .Q(n5732), .QN(n19286) );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(n3677), .CK(CLK), .RN(n20691), .Q(n5731), .QN(n19285) );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(n3676), .CK(CLK), .RN(n20740), .Q(n5810), .QN(n19284) );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(n3675), .CK(CLK), .RN(n20739), .Q(n5809), .QN(n19283) );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(n3674), .CK(CLK), .RN(n20714), .Q(n5808), .QN(n19282) );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(n3673), .CK(CLK), .RN(n20726), .Q(n5807), .QN(n19281) );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(n3672), .CK(CLK), .RN(n20706), .Q(n5806), .QN(n19280) );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(n3671), .CK(CLK), .RN(n20700), .Q(n5805), .QN(n19279) );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(n3670), .CK(CLK), .RN(n20694), .Q(n5804), .QN(n19278) );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(n3669), .CK(CLK), .RN(n20725), .Q(n5803), .QN(n19277) );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(n3668), .CK(CLK), .RN(n20720), .Q(n5802), 
        .QN(n19276) );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(n3667), .CK(CLK), .RN(n20721), .Q(n5801), 
        .QN(n19275) );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(n3666), .CK(CLK), .RN(n20740), .Q(n5800), 
        .QN(n19274) );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(n3665), .CK(CLK), .RN(n20708), .Q(n5799), 
        .QN(n19273) );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(n3664), .CK(CLK), .RN(n20725), .Q(n5798), 
        .QN(n19272) );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(n3663), .CK(CLK), .RN(n20718), .Q(n5797), 
        .QN(n19271) );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(n3662), .CK(CLK), .RN(n20722), .Q(n5796), 
        .QN(n19270) );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(n3661), .CK(CLK), .RN(n20701), .Q(n5795), 
        .QN(n19269) );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(n3660), .CK(CLK), .RN(n20707), .Q(n5794), 
        .QN(n19268) );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(n3659), .CK(CLK), .RN(n20711), .Q(n5793), 
        .QN(n19267) );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(n3658), .CK(CLK), .RN(n20726), .Q(n5791), .QN(n19682) );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(n3657), .CK(CLK), .RN(n20721), .Q(n5790), .QN(n19681) );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(n3656), .CK(CLK), .RN(n20732), .Q(n5789), .QN(n19680) );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(n3655), .CK(CLK), .RN(n20745), .Q(n5788), .QN(n19679) );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(n3654), .CK(CLK), .RN(n20732), .Q(n5890), .QN(n19678) );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(n3653), .CK(CLK), .RN(n20700), .Q(n5888), .QN(n19677) );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(n3652), .CK(CLK), .RN(n20732), .Q(n5887), .QN(n19676) );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(n3651), .CK(CLK), .RN(n20723), .Q(n5886), .QN(n19675) );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(n3650), .CK(CLK), .RN(n20692), .Q(n5889), .QN(n19674) );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(n3649), .CK(CLK), .RN(n20704), .Q(n5885), .QN(n19673) );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(n3648), .CK(CLK), .RN(n20717), .Q(n5884), .QN(n19672) );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(n3647), .CK(CLK), .RN(n20738), .Q(n5883), .QN(n19671) );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(n3646), .CK(CLK), .RN(n20744), .Q(n5787), .QN(n19670) );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(n3645), .CK(CLK), .RN(n20691), .Q(n5786), .QN(n19669) );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(n3644), .CK(CLK), .RN(n20714), .Q(n5785), .QN(n19668) );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(n3643), .CK(CLK), .RN(n20713), .Q(n5784), .QN(n19667) );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(n3642), .CK(CLK), .RN(n20714), .Q(n5783), .QN(n19666) );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(n3641), .CK(CLK), .RN(n20726), .Q(n5782), .QN(n19665) );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(n3640), .CK(CLK), .RN(n20733), .Q(n5781), .QN(n19664) );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(n3639), .CK(CLK), .RN(n20699), .Q(n5780), .QN(n19663) );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(n3638), .CK(CLK), .RN(n20706), .Q(n5779), .QN(n19662) );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(n3637), .CK(CLK), .RN(n20696), .Q(n5778), .QN(n19661) );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(n3636), .CK(CLK), .RN(n20716), .Q(n5777), 
        .QN(n19660) );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(n3635), .CK(CLK), .RN(n20713), .Q(n5776), 
        .QN(n19659) );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(n3634), .CK(CLK), .RN(n20730), .Q(n5775), 
        .QN(n19658) );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(n3633), .CK(CLK), .RN(n20717), .Q(n5774), 
        .QN(n19657) );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(n3632), .CK(CLK), .RN(n20730), .Q(n5773), 
        .QN(n19656) );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(n3631), .CK(CLK), .RN(n20718), .Q(n5772), 
        .QN(n19655) );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(n3630), .CK(CLK), .RN(n20711), .Q(n5771), 
        .QN(n19654) );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(n3629), .CK(CLK), .RN(n20728), .Q(n5770), 
        .QN(n19653) );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(n3628), .CK(CLK), .RN(n20729), .Q(n5769), 
        .QN(n19652) );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(n3627), .CK(CLK), .RN(n20713), .Q(n5768), 
        .QN(n19651) );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(n3626), .CK(CLK), .RN(n20694), .Q(
        n19202), .QN(n5509) );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(n3625), .CK(CLK), .RN(n20693), .Q(
        n19201), .QN(n5508) );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(n3624), .CK(CLK), .RN(n20705), .Q(
        n19200), .QN(n5507) );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(n3623), .CK(CLK), .RN(n20745), .Q(
        n19199), .QN(n5506) );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(n3622), .CK(CLK), .RN(n20744), .Q(
        n19198), .QN(n5505) );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(n3621), .CK(CLK), .RN(n20693), .Q(
        n19197), .QN(n5504) );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(n3620), .CK(CLK), .RN(n20701), .Q(
        n19196), .QN(n5503) );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(n3619), .CK(CLK), .RN(n20723), .Q(
        n19195), .QN(n5502) );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(n3618), .CK(CLK), .RN(n20744), .Q(
        n19194), .QN(n5475) );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(n3617), .CK(CLK), .RN(n20705), .Q(
        n19193), .QN(n5501) );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(n3616), .CK(CLK), .RN(n20717), .Q(
        n19192), .QN(n5500) );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(n3615), .CK(CLK), .RN(n20695), .Q(
        n19191), .QN(n5499) );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(n3614), .CK(CLK), .RN(n20744), .Q(
        n19190), .QN(n5498) );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(n3613), .CK(CLK), .RN(n20695), .Q(
        n19189), .QN(n5497) );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(n3612), .CK(CLK), .RN(n20736), .Q(
        n19188), .QN(n5496) );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(n3611), .CK(CLK), .RN(n20739), .Q(
        n19187), .QN(n5495) );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(n3610), .CK(CLK), .RN(n20714), .Q(
        n19186), .QN(n5494) );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(n3609), .CK(CLK), .RN(n20735), .Q(
        n19185), .QN(n5493) );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(n3608), .CK(CLK), .RN(n20693), .Q(
        n19184), .QN(n5492) );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(n3607), .CK(CLK), .RN(n20699), .Q(
        n19183), .QN(n5491) );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(n3606), .CK(CLK), .RN(n20739), .Q(
        n19182), .QN(n5490) );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(n3605), .CK(CLK), .RN(n20695), .Q(
        n19181), .QN(n5489) );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(n3604), .CK(CLK), .RN(n20707), .Q(n19180), .QN(n5488) );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(n3603), .CK(CLK), .RN(n20735), .Q(n19179), .QN(n5487) );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(n3602), .CK(CLK), .RN(n20722), .Q(n19178), .QN(n5486) );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(n3601), .CK(CLK), .RN(n20693), .Q(n19177), .QN(n5485) );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(n3600), .CK(CLK), .RN(n20700), .Q(n19176), .QN(n5484) );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(n3599), .CK(CLK), .RN(n20703), .Q(n19175), .QN(n5483) );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(n3598), .CK(CLK), .RN(n20695), .Q(n19174), .QN(n5482) );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(n3597), .CK(CLK), .RN(n20711), .Q(n19173), .QN(n5481) );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(n3596), .CK(CLK), .RN(n20730), .Q(n19172), .QN(n5480) );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(n3595), .CK(CLK), .RN(n20716), .Q(n19171), .QN(n5479) );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(n3594), .CK(CLK), .RN(n20719), .Q(n5006), .QN(n19746) );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(n3593), .CK(CLK), .RN(n20715), .Q(n5005), .QN(n19745) );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(n3592), .CK(CLK), .RN(n20698), .Q(n5004), .QN(n19744) );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(n3591), .CK(CLK), .RN(n20721), .Q(n5003), .QN(n19743) );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(n3590), .CK(CLK), .RN(n20708), .Q(n5014), .QN(n19742) );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(n3589), .CK(CLK), .RN(n20731), .Q(n5013), .QN(n19741) );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(n3588), .CK(CLK), .RN(n20732), .Q(n5012), .QN(n19740) );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(n3587), .CK(CLK), .RN(n20702), .Q(n5011), .QN(n19739) );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(n3586), .CK(CLK), .RN(n20738), .Q(n5010), .QN(n19738) );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(n3585), .CK(CLK), .RN(n20731), .Q(n5009), .QN(n19737) );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(n3584), .CK(CLK), .RN(n20703), .Q(n5008), .QN(n19736) );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(n3583), .CK(CLK), .RN(n20724), .Q(n5007), .QN(n19735) );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(n3582), .CK(CLK), .RN(n20715), .Q(n5002), .QN(n19734) );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(n3581), .CK(CLK), .RN(n20698), .Q(n5001), .QN(n19733) );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(n3580), .CK(CLK), .RN(n20703), .Q(n5151), .QN(n19732) );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(n3579), .CK(CLK), .RN(n20693), .Q(n5093), .QN(n19731) );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(n3578), .CK(CLK), .RN(n20728), .Q(n5092), .QN(n19730) );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(n3577), .CK(CLK), .RN(n20742), .Q(n5091), .QN(n19729) );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(n3576), .CK(CLK), .RN(n20693), .Q(n5090), .QN(n19728) );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(n3575), .CK(CLK), .RN(n20730), .Q(n5089), .QN(n19727) );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(n3574), .CK(CLK), .RN(n20702), .Q(n5088), .QN(n19726) );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(n3573), .CK(CLK), .RN(n20692), .Q(n5087), .QN(n19725) );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(n3572), .CK(CLK), .RN(n20710), .Q(n5086), 
        .QN(n19724) );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(n3571), .CK(CLK), .RN(n20720), .Q(n5085), 
        .QN(n19723) );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(n3570), .CK(CLK), .RN(n20734), .Q(n5084), 
        .QN(n19722) );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(n3569), .CK(CLK), .RN(n20726), .Q(n5083), 
        .QN(n19721) );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(n3568), .CK(CLK), .RN(n20711), .Q(n5082), 
        .QN(n19720) );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(n3567), .CK(CLK), .RN(n20738), .Q(n5081), 
        .QN(n19719) );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(n3566), .CK(CLK), .RN(n20743), .Q(n5080), 
        .QN(n19718) );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(n3565), .CK(CLK), .RN(n20728), .Q(n5079), 
        .QN(n19717) );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(n3564), .CK(CLK), .RN(n20743), .Q(n5078), 
        .QN(n19716) );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(n3563), .CK(CLK), .RN(n20743), .Q(n5077), 
        .QN(n19715) );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(n3562), .CK(CLK), .RN(n20735), .QN(
        n18874) );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(n3561), .CK(CLK), .RN(n20721), .QN(
        n18873) );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(n3560), .CK(CLK), .RN(n20705), .QN(
        n18872) );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(n3559), .CK(CLK), .RN(n20745), .QN(
        n18871) );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(n3558), .CK(CLK), .RN(n20732), .QN(
        n18882) );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(n3557), .CK(CLK), .RN(n20707), .QN(
        n18880) );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(n3556), .CK(CLK), .RN(n20702), .QN(
        n18879) );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(n3555), .CK(CLK), .RN(n20723), .QN(
        n18878) );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(n3554), .CK(CLK), .RN(n20738), .QN(
        n18881) );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(n3553), .CK(CLK), .RN(n20734), .QN(
        n18877) );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(n3552), .CK(CLK), .RN(n20719), .QN(
        n18876) );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(n3551), .CK(CLK), .RN(n20715), .QN(
        n18875) );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(n3550), .CK(CLK), .RN(n20744), .QN(
        n18870) );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(n3549), .CK(CLK), .RN(n20695), .QN(
        n18869) );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(n3548), .CK(CLK), .RN(n20698), .QN(
        n18868) );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(n3547), .CK(CLK), .RN(n20727), .QN(
        n18867) );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(n3546), .CK(CLK), .RN(n20733), .QN(
        n18866) );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(n3545), .CK(CLK), .RN(n20735), .QN(
        n18865) );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(n3544), .CK(CLK), .RN(n20702), .QN(
        n18864) );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(n3543), .CK(CLK), .RN(n20692), .QN(
        n18863) );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(n3542), .CK(CLK), .RN(n20698), .QN(
        n18862) );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(n3541), .CK(CLK), .RN(n20716), .QN(
        n18861) );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(n3540), .CK(CLK), .RN(n20720), .QN(
        n18860) );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(n3539), .CK(CLK), .RN(n20713), .QN(
        n18859) );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(n3538), .CK(CLK), .RN(n20727), .QN(
        n18858) );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(n3537), .CK(CLK), .RN(n20708), .QN(
        n18857) );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(n3536), .CK(CLK), .RN(n20703), .QN(
        n18856) );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(n3535), .CK(CLK), .RN(n20726), .QN(
        n18855) );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(n3534), .CK(CLK), .RN(n20711), .QN(
        n18854) );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(n3533), .CK(CLK), .RN(n20701), .QN(
        n18853) );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(n3532), .CK(CLK), .RN(n20707), .QN(
        n18852) );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(n3531), .CK(CLK), .RN(n20716), .QN(
        n18851) );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(n3530), .CK(CLK), .RN(n20726), .Q(n4996), .QN(n19416) );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(n3529), .CK(CLK), .RN(n20721), .Q(n4995), .QN(n19415) );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(n3528), .CK(CLK), .RN(n20731), .Q(n4994), .QN(n19426) );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(n3527), .CK(CLK), .RN(n20745), .Q(n4993), .QN(n19414) );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(n3526), .CK(CLK), .RN(n20735), .Q(n4992), .QN(n19413) );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(n3525), .CK(CLK), .RN(n20693), .Q(n4991), .QN(n19425) );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(n3524), .CK(CLK), .RN(n20709), .Q(n4990), .QN(n19412) );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(n3523), .CK(CLK), .RN(n20723), .Q(n4989), .QN(n19411) );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(n3522), .CK(CLK), .RN(n20738), .Q(n4988), .QN(n19424) );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(n3521), .CK(CLK), .RN(n20734), .Q(n4987), .QN(n19410) );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(n3520), .CK(CLK), .RN(n20717), .Q(n4986), .QN(n19409) );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(n3519), .CK(CLK), .RN(n20695), .Q(n4985), .QN(n19423) );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(n3518), .CK(CLK), .RN(n20744), .Q(n4984), .QN(n19408) );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(n3517), .CK(CLK), .RN(n20714), .Q(n4983), .QN(n19407) );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(n3516), .CK(CLK), .RN(n20699), .Q(n4982), .QN(n19422) );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(n3515), .CK(CLK), .RN(n20705), .Q(n4981), .QN(n19406) );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(n3514), .CK(CLK), .RN(n20692), .Q(n4980), .QN(n19405) );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(n3513), .CK(CLK), .RN(n20735), .Q(n4979), .QN(n19421) );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(n3512), .CK(CLK), .RN(n20702), .Q(n4978), .QN(n19404) );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(n3511), .CK(CLK), .RN(n20735), .Q(n4933), .QN(n19403) );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(n3510), .CK(CLK), .RN(n20739), .Q(n4932), .QN(n19420) );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(n3509), .CK(CLK), .RN(n20741), .Q(n4931), .QN(n19402) );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(n3508), .CK(CLK), .RN(n20741), .Q(n4930), 
        .QN(n19401) );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(n3507), .CK(CLK), .RN(n20713), .Q(n4929), 
        .QN(n19419) );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(n3506), .CK(CLK), .RN(n20723), .Q(n4928), 
        .QN(n19400) );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(n3505), .CK(CLK), .RN(n20735), .Q(n4927), 
        .QN(n19399) );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(n3504), .CK(CLK), .RN(n20702), .Q(n4926), 
        .QN(n19418) );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(n3503), .CK(CLK), .RN(n20726), .Q(n4925), 
        .QN(n19398) );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(n3502), .CK(CLK), .RN(n20742), .Q(n4924), 
        .QN(n19397) );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(n3501), .CK(CLK), .RN(n20705), .Q(n4923), 
        .QN(n19417) );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(n3500), .CK(CLK), .RN(n20715), .Q(n4922), 
        .QN(n19396) );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(n3499), .CK(CLK), .RN(n20716), .Q(n4921), 
        .QN(n19395) );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(n3498), .CK(CLK), .RN(n20694), .Q(n5076), .QN(n18946) );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(n3497), .CK(CLK), .RN(n20708), .Q(n5075), .QN(n18945) );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(n3496), .CK(CLK), .RN(n20729), .Q(n5074), .QN(n18944) );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(n3495), .CK(CLK), .RN(n20721), .Q(n5073), .QN(n18943) );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(n3494), .CK(CLK), .RN(n20717), .Q(n5471), .QN(n18942) );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(n3493), .CK(CLK), .RN(n20724), .Q(n5469), .QN(n18941) );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(n3492), .CK(CLK), .RN(n20708), .Q(n5467), .QN(n18940) );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(n3491), .CK(CLK), .RN(n20723), .Q(n5465), .QN(n18939) );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(n3490), .CK(CLK), .RN(n20731), .Q(n5463), .QN(n18938) );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(n3489), .CK(CLK), .RN(n20705), .Q(n5461), .QN(n18937) );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(n3488), .CK(CLK), .RN(n20703), .Q(n5459), .QN(n18936) );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(n3487), .CK(CLK), .RN(n20724), .Q(n5457), .QN(n18935) );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(n3486), .CK(CLK), .RN(n20700), .Q(n5072), .QN(n18934) );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(n3485), .CK(CLK), .RN(n20698), .Q(n5071), .QN(n18933) );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(n3484), .CK(CLK), .RN(n20698), .Q(n5359), .QN(n18932) );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(n3483), .CK(CLK), .RN(n20705), .Q(n5358), .QN(n18931) );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(n3482), .CK(CLK), .RN(n20719), .Q(n5357), .QN(n18930) );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(n3481), .CK(CLK), .RN(n20742), .Q(n5356), .QN(n18929) );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(n3480), .CK(CLK), .RN(n20722), .Q(n5355), .QN(n18928) );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(n3479), .CK(CLK), .RN(n20702), .Q(n5354), .QN(n18927) );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(n3478), .CK(CLK), .RN(n20706), .Q(n5353), .QN(n18926) );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(n3477), .CK(CLK), .RN(n20696), .Q(n5352), .QN(n18925) );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(n3476), .CK(CLK), .RN(n20715), .Q(n5351), 
        .QN(n18924) );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(n3475), .CK(CLK), .RN(n20720), .Q(n5350), 
        .QN(n18923) );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(n3474), .CK(CLK), .RN(n20728), .Q(n5349), 
        .QN(n18922) );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(n3473), .CK(CLK), .RN(n20717), .Q(n5348), 
        .QN(n18921) );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(n3472), .CK(CLK), .RN(n20697), .Q(n5347), 
        .QN(n18920) );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(n3471), .CK(CLK), .RN(n20726), .Q(n5346), 
        .QN(n18919) );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(n3470), .CK(CLK), .RN(n20743), .Q(n5345), 
        .QN(n18918) );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(n3469), .CK(CLK), .RN(n20711), .Q(n5344), 
        .QN(n18917) );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(n3468), .CK(CLK), .RN(n20707), .Q(n5343), 
        .QN(n18916) );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(n3467), .CK(CLK), .RN(n20705), .Q(n5342), 
        .QN(n18915) );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(n3466), .CK(CLK), .RN(n20726), .Q(n5383), .QN(n19714) );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(n3465), .CK(CLK), .RN(n20732), .Q(n5382), .QN(n19713) );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(n3464), .CK(CLK), .RN(n20696), .Q(n5381), .QN(n19712) );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(n3463), .CK(CLK), .RN(n20721), .Q(n5380), .QN(n19711) );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(n3462), .CK(CLK), .RN(n20708), .Q(n5447), .QN(n19710) );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(n3461), .CK(CLK), .RN(n20731), .Q(n5446), .QN(n19709) );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(n3460), .CK(CLK), .RN(n20702), .Q(n5445), .QN(n19708) );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(n3459), .CK(CLK), .RN(n20723), .Q(n5444), .QN(n19707) );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(n3458), .CK(CLK), .RN(n20738), .Q(n5443), .QN(n19706) );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(n3457), .CK(CLK), .RN(n20734), .Q(n5442), .QN(n19705) );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(n3456), .CK(CLK), .RN(n20719), .Q(n5441), .QN(n19704) );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(n3455), .CK(CLK), .RN(n20727), .Q(n5440), .QN(n19703) );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(n3454), .CK(CLK), .RN(n20700), .Q(n5379), .QN(n19702) );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(n3453), .CK(CLK), .RN(n20714), .Q(n5378), .QN(n19701) );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(n3452), .CK(CLK), .RN(n20703), .Q(n5377), .QN(n19700) );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(n3451), .CK(CLK), .RN(n20705), .Q(n5376), .QN(n19699) );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(n3450), .CK(CLK), .RN(n20704), .Q(n5375), .QN(n19698) );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(n3449), .CK(CLK), .RN(n20742), .Q(n5374), .QN(n19697) );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(n3448), .CK(CLK), .RN(n20722), .Q(n5373), .QN(n19696) );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(n3447), .CK(CLK), .RN(n20729), .Q(n5372), .QN(n19695) );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(n3446), .CK(CLK), .RN(n20697), .Q(n5371), .QN(n19694) );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(n3445), .CK(CLK), .RN(n20746), .Q(n5370), .QN(n19693) );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(n3444), .CK(CLK), .RN(n20710), .Q(n5369), 
        .QN(n19692) );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(n3443), .CK(CLK), .RN(n20720), .Q(n5368), 
        .QN(n19691) );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(n3442), .CK(CLK), .RN(n20723), .Q(n5367), 
        .QN(n19690) );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(n3441), .CK(CLK), .RN(n20708), .Q(n5366), 
        .QN(n19689) );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(n3440), .CK(CLK), .RN(n20697), .Q(n5365), 
        .QN(n19688) );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(n3439), .CK(CLK), .RN(n20738), .Q(n5364), 
        .QN(n19687) );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(n3438), .CK(CLK), .RN(n20712), .Q(n5363), 
        .QN(n19686) );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(n3437), .CK(CLK), .RN(n20728), .Q(n5362), 
        .QN(n19685) );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(n3436), .CK(CLK), .RN(n20713), .Q(n5361), 
        .QN(n19684) );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(n3435), .CK(CLK), .RN(n20713), .Q(n5360), 
        .QN(n19683) );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(n3434), .CK(CLK), .RN(n20719), .Q(n5341), .QN(n19331) );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(n3429), .CK(CLK), .RN(n20732), .Q(n5340), .QN(n19362) );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(n3424), .CK(CLK), .RN(n20698), .Q(n5339), .QN(n19354) );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(n3419), .CK(CLK), .RN(n20721), .Q(n5338), .QN(n19353) );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(n3414), .CK(CLK), .RN(n20708), .Q(n5337), .QN(n19361) );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(n3409), .CK(CLK), .RN(n20731), .Q(n5335), .QN(n19352) );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(n3404), .CK(CLK), .RN(n20701), .Q(n5205), .QN(n19351) );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(n3399), .CK(CLK), .RN(n20695), .Q(n5203), .QN(n19350) );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(n3394), .CK(CLK), .RN(n20731), .Q(n5201), .QN(n19360) );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(n3389), .CK(CLK), .RN(n20734), .Q(n5199), .QN(n19349) );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(n3384), .CK(CLK), .RN(n20696), .Q(n5197), .QN(n19348) );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(n3379), .CK(CLK), .RN(n20724), .Q(n5196), .QN(n19347) );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(n3374), .CK(CLK), .RN(n20715), .Q(n5195), .QN(n19346) );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(n3369), .CK(CLK), .RN(n20714), .Q(n5194), .QN(n19345) );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(n3364), .CK(CLK), .RN(n20703), .Q(n5193), .QN(n19344) );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(n3359), .CK(CLK), .RN(n20718), .Q(n5192), .QN(n19359) );
  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(n3354), .CK(CLK), .RN(n20728), .Q(n5191), .QN(n19343) );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(n3349), .CK(CLK), .RN(n20702), .Q(n5190), .QN(n19342) );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(n3344), .CK(CLK), .RN(n20743), .Q(n5189), .QN(n19341) );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(n3339), .CK(CLK), .RN(n20729), .Q(n5188), .QN(n19358) );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(n3334), .CK(CLK), .RN(n20724), .Q(n5187), .QN(n19340) );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(n3329), .CK(CLK), .RN(n20741), .Q(n5186), .QN(n19339) );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(n3324), .CK(CLK), .RN(n20710), .Q(n5185), 
        .QN(n19357) );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(n3319), .CK(CLK), .RN(n20719), .Q(n5184), 
        .QN(n19338) );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(n3314), .CK(CLK), .RN(n20723), .Q(n5183), 
        .QN(n19337) );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(n3309), .CK(CLK), .RN(n20691), .Q(n5182), 
        .QN(n19336) );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(n3304), .CK(CLK), .RN(n20700), .Q(n5181), 
        .QN(n19356) );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(n3299), .CK(CLK), .RN(n20700), .Q(n5180), 
        .QN(n19335) );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(n3294), .CK(CLK), .RN(n20718), .Q(n5179), 
        .QN(n19334) );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(n3289), .CK(CLK), .RN(n20711), .Q(n5178), 
        .QN(n19333) );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(n3284), .CK(CLK), .RN(n20713), .Q(n5177), 
        .QN(n19355) );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(n3279), .CK(CLK), .RN(n20738), .Q(n5176), 
        .QN(n19332) );
  NOR3_X2 U2161 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n2675), .ZN(n2673) );
  NOR3_X2 U3544 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n5707), .ZN(n5699) );
  NAND3_X1 U3618 ( .A1(n1149), .A2(n1150), .A3(n1151), .ZN(n1148) );
  NAND3_X1 U3619 ( .A1(n1149), .A2(n1150), .A3(n1188), .ZN(n1187) );
  NAND3_X1 U3620 ( .A1(n1149), .A2(n1150), .A3(n1225), .ZN(n1191) );
  NAND3_X1 U3621 ( .A1(n2645), .A2(n2646), .A3(ENABLE), .ZN(n1078) );
  XOR2_X1 U3622 ( .A(ADD_WR[4]), .B(ADD_RD2[4]), .Z(n2652) );
  XOR2_X1 U3623 ( .A(ADD_WR[3]), .B(ADD_RD2[3]), .Z(n2651) );
  XOR2_X1 U3624 ( .A(ADD_WR[2]), .B(ADD_RD2[2]), .Z(n2650) );
  XOR2_X1 U3625 ( .A(n2653), .B(ADD_WR[0]), .Z(n2648) );
  XOR2_X1 U3626 ( .A(n2654), .B(ADD_WR[1]), .Z(n2647) );
  NAND3_X1 U3627 ( .A1(n5684), .A2(n5722), .A3(ENABLE), .ZN(n2750) );
  XOR2_X1 U3628 ( .A(ADD_WR[4]), .B(ADD_RD1[4]), .Z(n5728) );
  XOR2_X1 U3629 ( .A(ADD_WR[3]), .B(ADD_RD1[3]), .Z(n5727) );
  XOR2_X1 U3630 ( .A(ADD_WR[2]), .B(ADD_RD1[2]), .Z(n5726) );
  XOR2_X1 U3631 ( .A(n5707), .B(ADD_WR[0]), .Z(n5724) );
  XOR2_X1 U3632 ( .A(n5718), .B(ADD_WR[1]), .Z(n5723) );
  NAND3_X1 U3633 ( .A1(n5722), .A2(n20746), .A3(ENABLE), .ZN(n2697) );
  NAND3_X1 U3634 ( .A1(n2646), .A2(n20746), .A3(ENABLE), .ZN(n1838) );
  TBUF_X1 \OUT2_tri[0]  ( .A(n3015), .EN(n3016), .Z(OUT2[0]) );
  TBUF_X1 \OUT2_tri[1]  ( .A(n3013), .EN(n3014), .Z(OUT2[1]) );
  TBUF_X1 \OUT2_tri[2]  ( .A(n3011), .EN(n3012), .Z(OUT2[2]) );
  TBUF_X1 \OUT2_tri[3]  ( .A(n3009), .EN(n3010), .Z(OUT2[3]) );
  TBUF_X1 \OUT2_tri[4]  ( .A(n3007), .EN(n3008), .Z(OUT2[4]) );
  TBUF_X1 \OUT2_tri[5]  ( .A(n3005), .EN(n3006), .Z(OUT2[5]) );
  TBUF_X1 \OUT2_tri[6]  ( .A(n3003), .EN(n3004), .Z(OUT2[6]) );
  TBUF_X1 \OUT2_tri[7]  ( .A(n3001), .EN(n3002), .Z(OUT2[7]) );
  TBUF_X1 \OUT2_tri[8]  ( .A(n2999), .EN(n3000), .Z(OUT2[8]) );
  TBUF_X1 \OUT2_tri[9]  ( .A(n2997), .EN(n2998), .Z(OUT2[9]) );
  TBUF_X1 \OUT2_tri[10]  ( .A(n2995), .EN(n2996), .Z(OUT2[10]) );
  TBUF_X1 \OUT2_tri[11]  ( .A(n2993), .EN(n2994), .Z(OUT2[11]) );
  TBUF_X1 \OUT2_tri[12]  ( .A(n2991), .EN(n2992), .Z(OUT2[12]) );
  TBUF_X1 \OUT2_tri[13]  ( .A(n2989), .EN(n2990), .Z(OUT2[13]) );
  TBUF_X1 \OUT2_tri[14]  ( .A(n2987), .EN(n2988), .Z(OUT2[14]) );
  TBUF_X1 \OUT2_tri[15]  ( .A(n2985), .EN(n2986), .Z(OUT2[15]) );
  TBUF_X1 \OUT2_tri[16]  ( .A(n2983), .EN(n2984), .Z(OUT2[16]) );
  TBUF_X1 \OUT2_tri[17]  ( .A(n2981), .EN(n2982), .Z(OUT2[17]) );
  TBUF_X1 \OUT2_tri[18]  ( .A(n2979), .EN(n2980), .Z(OUT2[18]) );
  TBUF_X1 \OUT2_tri[19]  ( .A(n2977), .EN(n2978), .Z(OUT2[19]) );
  TBUF_X1 \OUT2_tri[20]  ( .A(n2975), .EN(n2976), .Z(OUT2[20]) );
  TBUF_X1 \OUT2_tri[21]  ( .A(n2973), .EN(n2974), .Z(OUT2[21]) );
  TBUF_X1 \OUT2_tri[22]  ( .A(n2971), .EN(n2972), .Z(OUT2[22]) );
  TBUF_X1 \OUT2_tri[23]  ( .A(n2969), .EN(n2970), .Z(OUT2[23]) );
  TBUF_X1 \OUT2_tri[24]  ( .A(n2967), .EN(n2968), .Z(OUT2[24]) );
  TBUF_X1 \OUT2_tri[25]  ( .A(n2965), .EN(n2966), .Z(OUT2[25]) );
  TBUF_X1 \OUT2_tri[26]  ( .A(n2963), .EN(n2964), .Z(OUT2[26]) );
  TBUF_X1 \OUT2_tri[27]  ( .A(n2961), .EN(n2962), .Z(OUT2[27]) );
  TBUF_X1 \OUT2_tri[28]  ( .A(n2959), .EN(n2960), .Z(OUT2[28]) );
  TBUF_X1 \OUT2_tri[29]  ( .A(n2957), .EN(n2958), .Z(OUT2[29]) );
  TBUF_X1 \OUT2_tri[30]  ( .A(n2955), .EN(n2956), .Z(OUT2[30]) );
  TBUF_X1 \OUT2_tri[31]  ( .A(n2953), .EN(n2954), .Z(OUT2[31]) );
  DFFRS_X1 \OUT2_tri_enable_reg[31]  ( .D(n4459), .CK(CLK), .RN(n20683), .SN(
        n20688), .Q(n2954), .QN(n4458) );
  DFFRS_X1 \OUT2_tri_enable_reg[30]  ( .D(n4457), .CK(CLK), .RN(n20683), .SN(
        n20691), .Q(n2956), .QN(n4456) );
  DFFRS_X1 \OUT2_tri_enable_reg[29]  ( .D(n4455), .CK(CLK), .RN(n20683), .SN(
        n20690), .Q(n2958), .QN(n4454) );
  DFFRS_X1 \OUT2_tri_enable_reg[28]  ( .D(n4453), .CK(CLK), .RN(n20683), .SN(
        n20690), .Q(n2960), .QN(n4452) );
  DFFRS_X1 \OUT2_tri_enable_reg[27]  ( .D(n4451), .CK(CLK), .RN(n20683), .SN(
        n20690), .Q(n2962), .QN(n4450) );
  DFFRS_X1 \OUT2_tri_enable_reg[26]  ( .D(n4449), .CK(CLK), .RN(n20683), .SN(
        n20690), .Q(n2964), .QN(n4448) );
  DFFRS_X1 \OUT2_tri_enable_reg[25]  ( .D(n4447), .CK(CLK), .RN(n20683), .SN(
        n20690), .Q(n2966), .QN(n4446) );
  DFFRS_X1 \OUT2_tri_enable_reg[24]  ( .D(n4445), .CK(CLK), .RN(n20683), .SN(
        n20690), .Q(n2968), .QN(n4444) );
  DFFRS_X1 \OUT2_tri_enable_reg[23]  ( .D(n4443), .CK(CLK), .RN(n20683), .SN(
        n20690), .Q(n2970), .QN(n4442) );
  DFFRS_X1 \OUT2_tri_enable_reg[22]  ( .D(n4441), .CK(CLK), .RN(n20683), .SN(
        n20690), .Q(n2972), .QN(n4440) );
  DFFRS_X1 \OUT2_tri_enable_reg[21]  ( .D(n4439), .CK(CLK), .RN(n20683), .SN(
        n20690), .Q(n2974), .QN(n4438) );
  DFFRS_X1 \OUT2_tri_enable_reg[20]  ( .D(n4437), .CK(CLK), .RN(n20683), .SN(
        n20690), .Q(n2976), .QN(n4436) );
  DFFRS_X1 \OUT2_tri_enable_reg[19]  ( .D(n4435), .CK(CLK), .RN(n20684), .SN(
        n20690), .Q(n2978), .QN(n4434) );
  DFFRS_X1 \OUT2_tri_enable_reg[18]  ( .D(n4433), .CK(CLK), .RN(n20684), .SN(
        n20690), .Q(n2980), .QN(n4432) );
  DFFRS_X1 \OUT2_tri_enable_reg[17]  ( .D(n4431), .CK(CLK), .RN(n20684), .SN(
        n20690), .Q(n2982), .QN(n4430) );
  DFFRS_X1 \OUT2_tri_enable_reg[16]  ( .D(n4429), .CK(CLK), .RN(n20684), .SN(
        n20689), .Q(n2984), .QN(n4428) );
  DFFRS_X1 \OUT2_tri_enable_reg[15]  ( .D(n4427), .CK(CLK), .RN(n20684), .SN(
        n20689), .Q(n2986), .QN(n4426) );
  DFFRS_X1 \OUT2_tri_enable_reg[14]  ( .D(n4425), .CK(CLK), .RN(n20684), .SN(
        n20689), .Q(n2988), .QN(n4424) );
  DFFRS_X1 \OUT2_tri_enable_reg[13]  ( .D(n4423), .CK(CLK), .RN(n20684), .SN(
        n20689), .Q(n2990), .QN(n4422) );
  DFFRS_X1 \OUT2_tri_enable_reg[12]  ( .D(n4421), .CK(CLK), .RN(n20684), .SN(
        n20689), .Q(n2992), .QN(n4420) );
  DFFRS_X1 \OUT2_tri_enable_reg[11]  ( .D(n4419), .CK(CLK), .RN(n20684), .SN(
        n20689), .Q(n2994), .QN(n4418) );
  DFFRS_X1 \OUT2_tri_enable_reg[10]  ( .D(n4417), .CK(CLK), .RN(n20684), .SN(
        n20689), .Q(n2996), .QN(n4416) );
  DFFRS_X1 \OUT2_tri_enable_reg[9]  ( .D(n4415), .CK(CLK), .RN(n20684), .SN(
        n20689), .Q(n2998), .QN(n4414) );
  DFFRS_X1 \OUT2_tri_enable_reg[8]  ( .D(n4413), .CK(CLK), .RN(n20684), .SN(
        n20689), .Q(n3000), .QN(n4412) );
  DFFRS_X1 \OUT2_tri_enable_reg[7]  ( .D(n4411), .CK(CLK), .RN(n20685), .SN(
        n20689), .Q(n3002), .QN(n4410) );
  DFFRS_X1 \OUT2_tri_enable_reg[6]  ( .D(n4409), .CK(CLK), .RN(n20685), .SN(
        n20689), .Q(n3004), .QN(n4408) );
  DFFRS_X1 \OUT2_tri_enable_reg[5]  ( .D(n4407), .CK(CLK), .RN(n20685), .SN(
        n20689), .Q(n3006), .QN(n4406) );
  DFFRS_X1 \OUT2_tri_enable_reg[4]  ( .D(n4405), .CK(CLK), .RN(n20685), .SN(
        n20689), .Q(n3008), .QN(n4404) );
  DFFRS_X1 \OUT2_tri_enable_reg[3]  ( .D(n4403), .CK(CLK), .RN(n20685), .SN(
        n20688), .Q(n3010), .QN(n4402) );
  DFFRS_X1 \OUT2_tri_enable_reg[2]  ( .D(n4401), .CK(CLK), .RN(n20685), .SN(
        n20688), .Q(n3012), .QN(n4400) );
  DFFRS_X1 \OUT2_tri_enable_reg[1]  ( .D(n4399), .CK(CLK), .RN(n20685), .SN(
        n20688), .Q(n3014), .QN(n4398) );
  DFFRS_X1 \OUT2_tri_enable_reg[0]  ( .D(n4397), .CK(CLK), .RN(n20685), .SN(
        n20688), .Q(n3016), .QN(n4396) );
  DFFRS_X1 \OUT2_reg[31]  ( .D(n3433), .CK(CLK), .RN(n3430), .SN(n3431), .Q(
        n2953), .QN(n3432) );
  DFFRS_X1 \OUT2_reg[30]  ( .D(n3428), .CK(CLK), .RN(n3425), .SN(n3426), .Q(
        n2955), .QN(n3427) );
  DFFRS_X1 \OUT2_reg[29]  ( .D(n3423), .CK(CLK), .RN(n3420), .SN(n3421), .Q(
        n2957), .QN(n3422) );
  DFFRS_X1 \OUT2_reg[28]  ( .D(n3418), .CK(CLK), .RN(n3415), .SN(n3416), .Q(
        n2959), .QN(n3417) );
  DFFRS_X1 \OUT2_reg[27]  ( .D(n3413), .CK(CLK), .RN(n3410), .SN(n3411), .Q(
        n2961), .QN(n3412) );
  DFFRS_X1 \OUT2_reg[26]  ( .D(n3408), .CK(CLK), .RN(n3405), .SN(n3406), .Q(
        n2963), .QN(n3407) );
  DFFRS_X1 \OUT2_reg[25]  ( .D(n3403), .CK(CLK), .RN(n3400), .SN(n3401), .Q(
        n2965), .QN(n3402) );
  DFFRS_X1 \OUT2_reg[24]  ( .D(n3398), .CK(CLK), .RN(n3395), .SN(n3396), .Q(
        n2967), .QN(n3397) );
  DFFRS_X1 \OUT2_reg[23]  ( .D(n3393), .CK(CLK), .RN(n3390), .SN(n3391), .Q(
        n2969), .QN(n3392) );
  DFFRS_X1 \OUT2_reg[22]  ( .D(n3388), .CK(CLK), .RN(n3385), .SN(n3386), .Q(
        n2971), .QN(n3387) );
  DFFRS_X1 \OUT2_reg[21]  ( .D(n3383), .CK(CLK), .RN(n3380), .SN(n3381), .Q(
        n2973), .QN(n3382) );
  DFFRS_X1 \OUT2_reg[20]  ( .D(n3378), .CK(CLK), .RN(n3375), .SN(n3376), .Q(
        n2975), .QN(n3377) );
  DFFRS_X1 \OUT2_reg[19]  ( .D(n3373), .CK(CLK), .RN(n3370), .SN(n3371), .Q(
        n2977), .QN(n3372) );
  DFFRS_X1 \OUT2_reg[18]  ( .D(n3368), .CK(CLK), .RN(n3365), .SN(n3366), .Q(
        n2979), .QN(n3367) );
  DFFRS_X1 \OUT2_reg[17]  ( .D(n3363), .CK(CLK), .RN(n3360), .SN(n3361), .Q(
        n2981), .QN(n3362) );
  DFFRS_X1 \OUT2_reg[16]  ( .D(n3358), .CK(CLK), .RN(n3355), .SN(n3356), .Q(
        n2983), .QN(n3357) );
  DFFRS_X1 \OUT2_reg[15]  ( .D(n3353), .CK(CLK), .RN(n3350), .SN(n3351), .Q(
        n2985), .QN(n3352) );
  DFFRS_X1 \OUT2_reg[14]  ( .D(n3348), .CK(CLK), .RN(n3345), .SN(n3346), .Q(
        n2987), .QN(n3347) );
  DFFRS_X1 \OUT2_reg[13]  ( .D(n3343), .CK(CLK), .RN(n3340), .SN(n3341), .Q(
        n2989), .QN(n3342) );
  DFFRS_X1 \OUT2_reg[12]  ( .D(n3338), .CK(CLK), .RN(n3335), .SN(n3336), .Q(
        n2991), .QN(n3337) );
  DFFRS_X1 \OUT2_reg[11]  ( .D(n3333), .CK(CLK), .RN(n3330), .SN(n3331), .Q(
        n2993), .QN(n3332) );
  DFFRS_X1 \OUT2_reg[10]  ( .D(n3328), .CK(CLK), .RN(n3325), .SN(n3326), .Q(
        n2995), .QN(n3327) );
  DFFRS_X1 \OUT2_reg[9]  ( .D(n3323), .CK(CLK), .RN(n3320), .SN(n3321), .Q(
        n2997), .QN(n3322) );
  DFFRS_X1 \OUT2_reg[8]  ( .D(n3318), .CK(CLK), .RN(n3315), .SN(n3316), .Q(
        n2999), .QN(n3317) );
  DFFRS_X1 \OUT2_reg[7]  ( .D(n3313), .CK(CLK), .RN(n3310), .SN(n3311), .Q(
        n3001), .QN(n3312) );
  DFFRS_X1 \OUT2_reg[6]  ( .D(n3308), .CK(CLK), .RN(n3305), .SN(n3306), .Q(
        n3003), .QN(n3307) );
  DFFRS_X1 \OUT2_reg[5]  ( .D(n3303), .CK(CLK), .RN(n3300), .SN(n3301), .Q(
        n3005), .QN(n3302) );
  DFFRS_X1 \OUT2_reg[4]  ( .D(n3298), .CK(CLK), .RN(n3295), .SN(n3296), .Q(
        n3007), .QN(n3297) );
  DFFRS_X1 \OUT2_reg[3]  ( .D(n3293), .CK(CLK), .RN(n3290), .SN(n3291), .Q(
        n3009), .QN(n3292) );
  DFFRS_X1 \OUT2_reg[2]  ( .D(n3288), .CK(CLK), .RN(n3285), .SN(n3286), .Q(
        n3011), .QN(n3287) );
  DFFRS_X1 \OUT2_reg[1]  ( .D(n3283), .CK(CLK), .RN(n3280), .SN(n3281), .Q(
        n3013), .QN(n3282) );
  DFFRS_X1 \OUT2_reg[0]  ( .D(n3278), .CK(CLK), .RN(n3275), .SN(n3276), .Q(
        n3015), .QN(n3277) );
  DFFRS_X1 \OUT1_tri_enable_reg[31]  ( .D(n3270), .CK(CLK), .RN(n20680), .SN(
        n20688), .Q(n3018), .QN(n3269) );
  DFFRS_X1 \OUT1_tri_enable_reg[30]  ( .D(n3264), .CK(CLK), .RN(n20680), .SN(
        n20688), .Q(n3020), .QN(n3263) );
  DFFRS_X1 \OUT1_tri_enable_reg[29]  ( .D(n3258), .CK(CLK), .RN(n20680), .SN(
        n20688), .Q(n3022), .QN(n3257) );
  DFFRS_X1 \OUT1_tri_enable_reg[28]  ( .D(n3252), .CK(CLK), .RN(n20680), .SN(
        n20688), .Q(n3024), .QN(n3251) );
  DFFRS_X1 \OUT1_tri_enable_reg[27]  ( .D(n3246), .CK(CLK), .RN(n20680), .SN(
        n20688), .Q(n3026), .QN(n3245) );
  DFFRS_X1 \OUT1_tri_enable_reg[26]  ( .D(n3240), .CK(CLK), .RN(n20680), .SN(
        n20688), .Q(n3028), .QN(n3239) );
  DFFRS_X1 \OUT1_tri_enable_reg[25]  ( .D(n3234), .CK(CLK), .RN(n20680), .SN(
        n20688), .Q(n3030), .QN(n3233) );
  DFFRS_X1 \OUT1_tri_enable_reg[24]  ( .D(n3228), .CK(CLK), .RN(n20680), .SN(
        n20688), .Q(n3032), .QN(n3227) );
  DFFRS_X1 \OUT1_tri_enable_reg[23]  ( .D(n3222), .CK(CLK), .RN(n20680), .SN(
        n20687), .Q(n3034), .QN(n3221) );
  DFFRS_X1 \OUT1_tri_enable_reg[22]  ( .D(n3216), .CK(CLK), .RN(n20680), .SN(
        n20687), .Q(n3036), .QN(n3215) );
  DFFRS_X1 \OUT1_tri_enable_reg[21]  ( .D(n3210), .CK(CLK), .RN(n20680), .SN(
        n20687), .Q(n3038), .QN(n3209) );
  DFFRS_X1 \OUT1_tri_enable_reg[20]  ( .D(n3204), .CK(CLK), .RN(n20680), .SN(
        n20687), .Q(n3040), .QN(n3203) );
  DFFRS_X1 \OUT1_tri_enable_reg[19]  ( .D(n3198), .CK(CLK), .RN(n20681), .SN(
        n20687), .Q(n3042), .QN(n3197) );
  DFFRS_X1 \OUT1_tri_enable_reg[18]  ( .D(n3192), .CK(CLK), .RN(n20681), .SN(
        n20687), .Q(n3044), .QN(n3191) );
  DFFRS_X1 \OUT1_tri_enable_reg[17]  ( .D(n3186), .CK(CLK), .RN(n20681), .SN(
        n20687), .Q(n3046), .QN(n3185) );
  DFFRS_X1 \OUT1_tri_enable_reg[16]  ( .D(n3180), .CK(CLK), .RN(n20681), .SN(
        n20687), .Q(n3048), .QN(n3179) );
  DFFRS_X1 \OUT1_tri_enable_reg[15]  ( .D(n3174), .CK(CLK), .RN(n20681), .SN(
        n20687), .Q(n3050), .QN(n3173) );
  DFFRS_X1 \OUT1_tri_enable_reg[14]  ( .D(n3168), .CK(CLK), .RN(n20681), .SN(
        n20687), .Q(n3052), .QN(n3167) );
  DFFRS_X1 \OUT1_tri_enable_reg[13]  ( .D(n3162), .CK(CLK), .RN(n20681), .SN(
        n20687), .Q(n3054), .QN(n3161) );
  DFFRS_X1 \OUT1_tri_enable_reg[12]  ( .D(n3156), .CK(CLK), .RN(n20681), .SN(
        n20687), .Q(n3056), .QN(n3155) );
  DFFRS_X1 \OUT1_tri_enable_reg[11]  ( .D(n3150), .CK(CLK), .RN(n20681), .SN(
        n20687), .Q(n3058), .QN(n3149) );
  DFFRS_X1 \OUT1_tri_enable_reg[10]  ( .D(n3144), .CK(CLK), .RN(n20681), .SN(
        n20686), .Q(n3060), .QN(n3143) );
  DFFRS_X1 \OUT1_tri_enable_reg[9]  ( .D(n3138), .CK(CLK), .RN(n20681), .SN(
        n20686), .Q(n3062), .QN(n3137) );
  DFFRS_X1 \OUT1_tri_enable_reg[8]  ( .D(n3132), .CK(CLK), .RN(n20681), .SN(
        n20686), .Q(n3064), .QN(n3131) );
  DFFRS_X1 \OUT1_tri_enable_reg[7]  ( .D(n3126), .CK(CLK), .RN(n20682), .SN(
        n20686), .Q(n3066), .QN(n3125) );
  DFFRS_X1 \OUT1_tri_enable_reg[6]  ( .D(n3120), .CK(CLK), .RN(n20682), .SN(
        n20686), .Q(n3068), .QN(n3119) );
  DFFRS_X1 \OUT1_tri_enable_reg[5]  ( .D(n3114), .CK(CLK), .RN(n20682), .SN(
        n20686), .Q(n3070), .QN(n3113) );
  DFFRS_X1 \OUT1_tri_enable_reg[4]  ( .D(n3108), .CK(CLK), .RN(n20682), .SN(
        n20686), .Q(n3072), .QN(n3107) );
  DFFRS_X1 \OUT1_tri_enable_reg[3]  ( .D(n3102), .CK(CLK), .RN(n20682), .SN(
        n20686), .Q(n3074), .QN(n3101) );
  DFFRS_X1 \OUT1_tri_enable_reg[2]  ( .D(n3096), .CK(CLK), .RN(n20682), .SN(
        n20686), .Q(n3076), .QN(n3095) );
  DFFRS_X1 \OUT1_tri_enable_reg[1]  ( .D(n3090), .CK(CLK), .RN(n20682), .SN(
        n20686), .Q(n3078), .QN(n3089) );
  DFFRS_X1 \OUT1_tri_enable_reg[0]  ( .D(n3084), .CK(CLK), .RN(n20682), .SN(
        n20686), .Q(n3080), .QN(n3083) );
  DFFRS_X1 \OUT1_reg[30]  ( .D(n3268), .CK(CLK), .RN(n3265), .SN(n3266), .Q(
        n3019), .QN(n3267) );
  DFFRS_X1 \OUT1_reg[27]  ( .D(n3250), .CK(CLK), .RN(n3247), .SN(n3248), .Q(
        n3025), .QN(n3249) );
  DFFRS_X1 \OUT1_reg[23]  ( .D(n3226), .CK(CLK), .RN(n3223), .SN(n3224), .Q(
        n3033), .QN(n3225) );
  DFFRS_X1 \OUT1_reg[16]  ( .D(n3184), .CK(CLK), .RN(n3181), .SN(n3182), .Q(
        n3047), .QN(n3183) );
  DFFRS_X1 \OUT1_reg[12]  ( .D(n3160), .CK(CLK), .RN(n3157), .SN(n3158), .Q(
        n3055), .QN(n3159) );
  DFFRS_X1 \OUT1_reg[9]  ( .D(n3142), .CK(CLK), .RN(n3139), .SN(n3140), .Q(
        n3061), .QN(n3141) );
  DFFRS_X1 \OUT1_reg[5]  ( .D(n3118), .CK(CLK), .RN(n3115), .SN(n3116), .Q(
        n3069), .QN(n3117) );
  DFFRS_X1 \OUT1_reg[1]  ( .D(n3094), .CK(CLK), .RN(n3091), .SN(n3092), .Q(
        n3077), .QN(n3093) );
  DFFRS_X1 \OUT1_reg[31]  ( .D(n3274), .CK(CLK), .RN(n3271), .SN(n3272), .Q(
        n3017), .QN(n3273) );
  DFFRS_X1 \OUT1_reg[29]  ( .D(n3262), .CK(CLK), .RN(n3259), .SN(n3260), .Q(
        n3021), .QN(n3261) );
  DFFRS_X1 \OUT1_reg[28]  ( .D(n3256), .CK(CLK), .RN(n3253), .SN(n3254), .Q(
        n3023), .QN(n3255) );
  DFFRS_X1 \OUT1_reg[26]  ( .D(n3244), .CK(CLK), .RN(n3241), .SN(n3242), .Q(
        n3027), .QN(n3243) );
  DFFRS_X1 \OUT1_reg[25]  ( .D(n3238), .CK(CLK), .RN(n3235), .SN(n3236), .Q(
        n3029), .QN(n3237) );
  DFFRS_X1 \OUT1_reg[24]  ( .D(n3232), .CK(CLK), .RN(n3229), .SN(n3230), .Q(
        n3031), .QN(n3231) );
  DFFRS_X1 \OUT1_reg[22]  ( .D(n3220), .CK(CLK), .RN(n3217), .SN(n3218), .Q(
        n3035), .QN(n3219) );
  DFFRS_X1 \OUT1_reg[21]  ( .D(n3214), .CK(CLK), .RN(n3211), .SN(n3212), .Q(
        n3037), .QN(n3213) );
  DFFRS_X1 \OUT1_reg[20]  ( .D(n3208), .CK(CLK), .RN(n3205), .SN(n3206), .Q(
        n3039), .QN(n3207) );
  DFFRS_X1 \OUT1_reg[19]  ( .D(n3202), .CK(CLK), .RN(n3199), .SN(n3200), .Q(
        n3041), .QN(n3201) );
  DFFRS_X1 \OUT1_reg[18]  ( .D(n3196), .CK(CLK), .RN(n3193), .SN(n3194), .Q(
        n3043), .QN(n3195) );
  DFFRS_X1 \OUT1_reg[17]  ( .D(n3190), .CK(CLK), .RN(n3187), .SN(n3188), .Q(
        n3045), .QN(n3189) );
  DFFRS_X1 \OUT1_reg[15]  ( .D(n3178), .CK(CLK), .RN(n3175), .SN(n3176), .Q(
        n3049), .QN(n3177) );
  DFFRS_X1 \OUT1_reg[14]  ( .D(n3172), .CK(CLK), .RN(n3169), .SN(n3170), .Q(
        n3051), .QN(n3171) );
  DFFRS_X1 \OUT1_reg[13]  ( .D(n3166), .CK(CLK), .RN(n3163), .SN(n3164), .Q(
        n3053), .QN(n3165) );
  DFFRS_X1 \OUT1_reg[11]  ( .D(n3154), .CK(CLK), .RN(n3151), .SN(n3152), .Q(
        n3057), .QN(n3153) );
  DFFRS_X1 \OUT1_reg[10]  ( .D(n3148), .CK(CLK), .RN(n3145), .SN(n3146), .Q(
        n3059), .QN(n3147) );
  DFFRS_X1 \OUT1_reg[8]  ( .D(n3136), .CK(CLK), .RN(n3133), .SN(n3134), .Q(
        n3063), .QN(n3135) );
  DFFRS_X1 \OUT1_reg[7]  ( .D(n3130), .CK(CLK), .RN(n3127), .SN(n3128), .Q(
        n3065), .QN(n3129) );
  DFFRS_X1 \OUT1_reg[6]  ( .D(n3124), .CK(CLK), .RN(n3121), .SN(n3122), .Q(
        n3067), .QN(n3123) );
  DFFRS_X1 \OUT1_reg[4]  ( .D(n3112), .CK(CLK), .RN(n3109), .SN(n3110), .Q(
        n3071), .QN(n3111) );
  DFFRS_X1 \OUT1_reg[3]  ( .D(n3106), .CK(CLK), .RN(n3103), .SN(n3104), .Q(
        n3073), .QN(n3105) );
  DFFRS_X1 \OUT1_reg[2]  ( .D(n3100), .CK(CLK), .RN(n3097), .SN(n3098), .Q(
        n3075), .QN(n3099) );
  DFFRS_X1 \OUT1_reg[0]  ( .D(n3088), .CK(CLK), .RN(n3085), .SN(n3086), .Q(
        n3079), .QN(n3087) );
  TBUF_X1 \OUT1_tri[1]  ( .A(n3077), .EN(n3078), .Z(OUT1[1]) );
  TBUF_X1 \OUT1_tri[5]  ( .A(n3069), .EN(n3070), .Z(OUT1[5]) );
  TBUF_X1 \OUT1_tri[9]  ( .A(n3061), .EN(n3062), .Z(OUT1[9]) );
  TBUF_X1 \OUT1_tri[12]  ( .A(n3055), .EN(n3056), .Z(OUT1[12]) );
  TBUF_X1 \OUT1_tri[16]  ( .A(n3047), .EN(n3048), .Z(OUT1[16]) );
  TBUF_X1 \OUT1_tri[23]  ( .A(n3033), .EN(n3034), .Z(OUT1[23]) );
  TBUF_X1 \OUT1_tri[27]  ( .A(n3025), .EN(n3026), .Z(OUT1[27]) );
  TBUF_X1 \OUT1_tri[30]  ( .A(n3019), .EN(n3020), .Z(OUT1[30]) );
  TBUF_X1 \OUT1_tri[2]  ( .A(n3075), .EN(n3076), .Z(OUT1[2]) );
  TBUF_X1 \OUT1_tri[4]  ( .A(n3071), .EN(n3072), .Z(OUT1[4]) );
  TBUF_X1 \OUT1_tri[8]  ( .A(n3063), .EN(n3064), .Z(OUT1[8]) );
  TBUF_X1 \OUT1_tri[11]  ( .A(n3057), .EN(n3058), .Z(OUT1[11]) );
  TBUF_X1 \OUT1_tri[15]  ( .A(n3049), .EN(n3050), .Z(OUT1[15]) );
  TBUF_X1 \OUT1_tri[19]  ( .A(n3041), .EN(n3042), .Z(OUT1[19]) );
  TBUF_X1 \OUT1_tri[22]  ( .A(n3035), .EN(n3036), .Z(OUT1[22]) );
  TBUF_X1 \OUT1_tri[26]  ( .A(n3027), .EN(n3028), .Z(OUT1[26]) );
  TBUF_X1 \OUT1_tri[3]  ( .A(n3073), .EN(n3074), .Z(OUT1[3]) );
  TBUF_X1 \OUT1_tri[7]  ( .A(n3065), .EN(n3066), .Z(OUT1[7]) );
  TBUF_X1 \OUT1_tri[10]  ( .A(n3059), .EN(n3060), .Z(OUT1[10]) );
  TBUF_X1 \OUT1_tri[14]  ( .A(n3051), .EN(n3052), .Z(OUT1[14]) );
  TBUF_X1 \OUT1_tri[18]  ( .A(n3043), .EN(n3044), .Z(OUT1[18]) );
  TBUF_X1 \OUT1_tri[21]  ( .A(n3037), .EN(n3038), .Z(OUT1[21]) );
  TBUF_X1 \OUT1_tri[25]  ( .A(n3029), .EN(n3030), .Z(OUT1[25]) );
  TBUF_X1 \OUT1_tri[29]  ( .A(n3021), .EN(n3022), .Z(OUT1[29]) );
  TBUF_X1 \OUT1_tri[0]  ( .A(n3079), .EN(n3080), .Z(OUT1[0]) );
  TBUF_X1 \OUT1_tri[6]  ( .A(n3067), .EN(n3068), .Z(OUT1[6]) );
  TBUF_X1 \OUT1_tri[13]  ( .A(n3053), .EN(n3054), .Z(OUT1[13]) );
  TBUF_X1 \OUT1_tri[17]  ( .A(n3045), .EN(n3046), .Z(OUT1[17]) );
  TBUF_X1 \OUT1_tri[20]  ( .A(n3039), .EN(n3040), .Z(OUT1[20]) );
  TBUF_X1 \OUT1_tri[24]  ( .A(n3031), .EN(n3032), .Z(OUT1[24]) );
  TBUF_X1 \OUT1_tri[28]  ( .A(n3023), .EN(n3024), .Z(OUT1[28]) );
  TBUF_X1 \OUT1_tri[31]  ( .A(n3017), .EN(n3018), .Z(OUT1[31]) );
  NOR2_X1 U3 ( .A1(n5718), .A2(ADD_RD1[2]), .ZN(n5696) );
  NOR3_X1 U4 ( .A1(n2653), .A2(ADD_RD2[4]), .A3(n2675), .ZN(n2665) );
  NOR2_X1 U5 ( .A1(n2689), .A2(ADD_RD2[1]), .ZN(n2669) );
  NOR2_X1 U6 ( .A1(n2654), .A2(ADD_RD2[2]), .ZN(n2666) );
  NOR3_X1 U7 ( .A1(n5707), .A2(ADD_RD1[4]), .A3(n5710), .ZN(n5695) );
  NOR2_X1 U8 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n5703) );
  NOR2_X1 U9 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n2674) );
  NOR2_X1 U10 ( .A1(n1727), .A2(ADD_WR[2]), .ZN(n1151) );
  NOR2_X1 U11 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .ZN(n1146) );
  NOR2_X1 U12 ( .A1(n1796), .A2(n1727), .ZN(n1225) );
  NOR2_X1 U13 ( .A1(n1796), .A2(ADD_WR[1]), .ZN(n1188) );
  AND2_X1 U14 ( .A1(n1151), .A2(n1145), .ZN(n18850) );
  BUF_X1 U15 ( .A(n20402), .Z(n19809) );
  BUF_X1 U16 ( .A(n20402), .Z(n19810) );
  BUF_X1 U17 ( .A(n20401), .Z(n19811) );
  BUF_X1 U18 ( .A(n20374), .Z(n19800) );
  BUF_X1 U19 ( .A(n20374), .Z(n19801) );
  BUF_X1 U20 ( .A(n20446), .Z(n19824) );
  BUF_X1 U21 ( .A(n20446), .Z(n19825) );
  BUF_X1 U22 ( .A(n20464), .Z(n19830) );
  BUF_X1 U23 ( .A(n20464), .Z(n19831) );
  BUF_X1 U24 ( .A(n20514), .Z(n19848) );
  BUF_X1 U25 ( .A(n20514), .Z(n19849) );
  BUF_X1 U26 ( .A(n20480), .Z(n19836) );
  BUF_X1 U27 ( .A(n20480), .Z(n19837) );
  BUF_X1 U28 ( .A(n20496), .Z(n19842) );
  BUF_X1 U29 ( .A(n20496), .Z(n19843) );
  BUF_X1 U30 ( .A(n20506), .Z(n19845) );
  BUF_X1 U31 ( .A(n20506), .Z(n19846) );
  BUF_X1 U32 ( .A(n20523), .Z(n19851) );
  BUF_X1 U33 ( .A(n20523), .Z(n19852) );
  BUF_X1 U34 ( .A(n20464), .Z(n19832) );
  BUF_X1 U35 ( .A(n20514), .Z(n19850) );
  BUF_X1 U36 ( .A(n20505), .Z(n19847) );
  BUF_X1 U37 ( .A(n20524), .Z(n19853) );
  BUF_X1 U38 ( .A(n20419), .Z(n19815) );
  BUF_X1 U39 ( .A(n20419), .Z(n19816) );
  BUF_X1 U40 ( .A(n20455), .Z(n19827) );
  BUF_X1 U41 ( .A(n20455), .Z(n19828) );
  BUF_X1 U42 ( .A(n20320), .Z(n19782) );
  BUF_X1 U43 ( .A(n20320), .Z(n19783) );
  BUF_X1 U44 ( .A(n20329), .Z(n19785) );
  BUF_X1 U45 ( .A(n20329), .Z(n19786) );
  BUF_X1 U46 ( .A(n20339), .Z(n19788) );
  BUF_X1 U47 ( .A(n20339), .Z(n19789) );
  BUF_X1 U48 ( .A(n20347), .Z(n19791) );
  BUF_X1 U49 ( .A(n20347), .Z(n19792) );
  BUF_X1 U50 ( .A(n20357), .Z(n19794) );
  BUF_X1 U51 ( .A(n20357), .Z(n19795) );
  BUF_X1 U52 ( .A(n20365), .Z(n19797) );
  BUF_X1 U53 ( .A(n20365), .Z(n19798) );
  BUF_X1 U54 ( .A(n20383), .Z(n19803) );
  BUF_X1 U55 ( .A(n20383), .Z(n19804) );
  BUF_X1 U56 ( .A(n20392), .Z(n19806) );
  BUF_X1 U57 ( .A(n20392), .Z(n19807) );
  BUF_X1 U58 ( .A(n20410), .Z(n19812) );
  BUF_X1 U59 ( .A(n20410), .Z(n19813) );
  BUF_X1 U60 ( .A(n20428), .Z(n19818) );
  BUF_X1 U61 ( .A(n20428), .Z(n19819) );
  BUF_X1 U62 ( .A(n20437), .Z(n19821) );
  BUF_X1 U63 ( .A(n20437), .Z(n19822) );
  BUF_X1 U64 ( .A(n20374), .Z(n19802) );
  BUF_X1 U65 ( .A(n20419), .Z(n19817) );
  BUF_X1 U66 ( .A(n20446), .Z(n19826) );
  BUF_X1 U67 ( .A(n20455), .Z(n19829) );
  BUF_X1 U68 ( .A(n20321), .Z(n19784) );
  BUF_X1 U69 ( .A(n20330), .Z(n19787) );
  BUF_X1 U70 ( .A(n20338), .Z(n19790) );
  BUF_X1 U71 ( .A(n20348), .Z(n19793) );
  BUF_X1 U72 ( .A(n20356), .Z(n19796) );
  BUF_X1 U73 ( .A(n20366), .Z(n19799) );
  BUF_X1 U74 ( .A(n20384), .Z(n19805) );
  BUF_X1 U75 ( .A(n20393), .Z(n19808) );
  BUF_X1 U76 ( .A(n20411), .Z(n19814) );
  BUF_X1 U77 ( .A(n20429), .Z(n19820) );
  BUF_X1 U78 ( .A(n20438), .Z(n19823) );
  BUF_X1 U79 ( .A(n20481), .Z(n19838) );
  BUF_X1 U80 ( .A(n20497), .Z(n19844) );
  INV_X1 U81 ( .A(n20546), .ZN(n20536) );
  INV_X1 U82 ( .A(n20546), .ZN(n20537) );
  BUF_X1 U83 ( .A(n1367), .Z(n19839) );
  BUF_X1 U84 ( .A(n1367), .Z(n19840) );
  BUF_X1 U85 ( .A(n1186), .Z(n19863) );
  BUF_X1 U86 ( .A(n1186), .Z(n19864) );
  BUF_X1 U87 ( .A(n1192), .Z(n19857) );
  BUF_X1 U88 ( .A(n1192), .Z(n19858) );
  BUF_X1 U89 ( .A(n1403), .Z(n19833) );
  BUF_X1 U90 ( .A(n1403), .Z(n19834) );
  INV_X1 U91 ( .A(n20560), .ZN(n20551) );
  INV_X1 U92 ( .A(n20560), .ZN(n20550) );
  BUF_X1 U93 ( .A(n1367), .Z(n19841) );
  BUF_X1 U94 ( .A(n1186), .Z(n19865) );
  BUF_X1 U95 ( .A(n1192), .Z(n19859) );
  BUF_X1 U96 ( .A(n1403), .Z(n19835) );
  BUF_X1 U97 ( .A(n2695), .Z(n19780) );
  BUF_X1 U98 ( .A(n2695), .Z(n19779) );
  BUF_X1 U99 ( .A(n1189), .Z(n19860) );
  BUF_X1 U100 ( .A(n1189), .Z(n19861) );
  BUF_X1 U101 ( .A(n1227), .Z(n19854) );
  BUF_X1 U102 ( .A(n1227), .Z(n19855) );
  BUF_X1 U103 ( .A(n2695), .Z(n19781) );
  INV_X1 U104 ( .A(n20679), .ZN(n20670) );
  INV_X1 U105 ( .A(n20679), .ZN(n20669) );
  BUF_X1 U106 ( .A(n2693), .Z(n20104) );
  BUF_X1 U107 ( .A(n1834), .Z(n20317) );
  BUF_X1 U108 ( .A(n2693), .Z(n20105) );
  BUF_X1 U109 ( .A(n1834), .Z(n20318) );
  BUF_X1 U110 ( .A(n2693), .Z(n20106) );
  BUF_X1 U111 ( .A(n1834), .Z(n20319) );
  INV_X1 U112 ( .A(n2712), .ZN(n20073) );
  INV_X1 U113 ( .A(n2712), .ZN(n20074) );
  AND2_X1 U114 ( .A1(n2687), .A2(n2667), .ZN(n1882) );
  INV_X1 U115 ( .A(n1848), .ZN(n20298) );
  INV_X1 U116 ( .A(n1865), .ZN(n20227) );
  INV_X1 U117 ( .A(n2723), .ZN(n20016) );
  INV_X1 U118 ( .A(n2724), .ZN(n20024) );
  INV_X1 U119 ( .A(n1860), .ZN(n20259) );
  INV_X1 U120 ( .A(n1875), .ZN(n20211) );
  INV_X1 U121 ( .A(n1892), .ZN(n20131) );
  INV_X1 U122 ( .A(n1878), .ZN(n20187) );
  INV_X1 U123 ( .A(n1891), .ZN(n20123) );
  INV_X1 U124 ( .A(n1866), .ZN(n20235) );
  INV_X1 U125 ( .A(n1877), .ZN(n20179) );
  INV_X1 U126 ( .A(n1885), .ZN(n20155) );
  INV_X1 U127 ( .A(n1886), .ZN(n20163) );
  INV_X1 U128 ( .A(n2732), .ZN(n20000) );
  INV_X1 U129 ( .A(n2744), .ZN(n19952) );
  INV_X1 U130 ( .A(n2749), .ZN(n19921) );
  INV_X1 U131 ( .A(n2748), .ZN(n19913) );
  INV_X1 U132 ( .A(n2749), .ZN(n19920) );
  INV_X1 U133 ( .A(n2748), .ZN(n19912) );
  INV_X1 U134 ( .A(n2734), .ZN(n19968) );
  INV_X1 U135 ( .A(n2735), .ZN(n19976) );
  INV_X1 U136 ( .A(n2743), .ZN(n19945) );
  INV_X1 U137 ( .A(n2743), .ZN(n19944) );
  INV_X1 U138 ( .A(n2733), .ZN(n20008) );
  INV_X1 U139 ( .A(n1876), .ZN(n20219) );
  INV_X1 U140 ( .A(n1876), .ZN(n20220) );
  INV_X1 U141 ( .A(n2718), .ZN(n20049) );
  BUF_X1 U142 ( .A(n20287), .Z(n20288) );
  BUF_X1 U143 ( .A(n20287), .Z(n20289) );
  BUF_X1 U144 ( .A(n20306), .Z(n20307) );
  BUF_X1 U145 ( .A(n20306), .Z(n20308) );
  BUF_X1 U146 ( .A(n18850), .Z(n20546) );
  BUF_X1 U147 ( .A(n20091), .Z(n20092) );
  BUF_X1 U148 ( .A(n20091), .Z(n20093) );
  BUF_X1 U149 ( .A(n20040), .Z(n20041) );
  BUF_X1 U150 ( .A(n20040), .Z(n20042) );
  BUF_X1 U151 ( .A(n20084), .Z(n20085) );
  BUF_X1 U152 ( .A(n20084), .Z(n20086) );
  BUF_X1 U153 ( .A(n20287), .Z(n20290) );
  BUF_X1 U154 ( .A(n1854), .Z(n20291) );
  BUF_X1 U155 ( .A(n1854), .Z(n20292) );
  BUF_X1 U156 ( .A(n1854), .Z(n20293) );
  BUF_X1 U157 ( .A(n20306), .Z(n20309) );
  BUF_X1 U158 ( .A(n1849), .Z(n20310) );
  BUF_X1 U159 ( .A(n1849), .Z(n20311) );
  BUF_X1 U160 ( .A(n1849), .Z(n20312) );
  BUF_X1 U161 ( .A(n20091), .Z(n20094) );
  BUF_X1 U162 ( .A(n2707), .Z(n20095) );
  BUF_X1 U163 ( .A(n2707), .Z(n20097) );
  BUF_X1 U164 ( .A(n2707), .Z(n20096) );
  BUF_X1 U165 ( .A(n20040), .Z(n20043) );
  BUF_X1 U166 ( .A(n2727), .Z(n20044) );
  BUF_X1 U167 ( .A(n2727), .Z(n20046) );
  BUF_X1 U168 ( .A(n2727), .Z(n20045) );
  BUF_X1 U169 ( .A(n20084), .Z(n20087) );
  BUF_X1 U170 ( .A(n2716), .Z(n20088) );
  BUF_X1 U171 ( .A(n2716), .Z(n20090) );
  BUF_X1 U172 ( .A(n2716), .Z(n20089) );
  INV_X1 U173 ( .A(n20665), .ZN(n20657) );
  INV_X1 U174 ( .A(n20665), .ZN(n20658) );
  BUF_X1 U175 ( .A(n1189), .Z(n19862) );
  BUF_X1 U176 ( .A(n1227), .Z(n19856) );
  INV_X1 U177 ( .A(n1554), .ZN(n20401) );
  INV_X1 U178 ( .A(n1554), .ZN(n20402) );
  BUF_X1 U179 ( .A(n20549), .Z(n20560) );
  BUF_X1 U180 ( .A(n20549), .Z(n20559) );
  BUF_X1 U181 ( .A(n20549), .Z(n20558) );
  BUF_X1 U182 ( .A(n20548), .Z(n20557) );
  BUF_X1 U183 ( .A(n20548), .Z(n20556) );
  BUF_X1 U184 ( .A(n20548), .Z(n20555) );
  BUF_X1 U185 ( .A(n20547), .Z(n20554) );
  BUF_X1 U186 ( .A(n20547), .Z(n20553) );
  BUF_X1 U187 ( .A(n20547), .Z(n20552) );
  BUF_X1 U188 ( .A(n20540), .Z(n20545) );
  BUF_X1 U189 ( .A(n20541), .Z(n20544) );
  BUF_X1 U190 ( .A(n18850), .Z(n20543) );
  BUF_X1 U191 ( .A(n18850), .Z(n20542) );
  BUF_X1 U192 ( .A(n18850), .Z(n20541) );
  BUF_X1 U193 ( .A(n18850), .Z(n20540) );
  BUF_X1 U194 ( .A(n18850), .Z(n20539) );
  BUF_X1 U195 ( .A(n18850), .Z(n20538) );
  INV_X1 U196 ( .A(n19892), .ZN(n1192) );
  INV_X1 U197 ( .A(n19895), .ZN(n1186) );
  INV_X1 U198 ( .A(n20479), .ZN(n1403) );
  INV_X1 U199 ( .A(n20495), .ZN(n1367) );
  BUF_X1 U200 ( .A(n18776), .Z(n20681) );
  BUF_X1 U201 ( .A(n18776), .Z(n20680) );
  BUF_X1 U202 ( .A(n18773), .Z(n20684) );
  BUF_X1 U203 ( .A(n18773), .Z(n20683) );
  BUF_X1 U204 ( .A(n18776), .Z(n20682) );
  BUF_X1 U205 ( .A(n18773), .Z(n20685) );
  NOR2_X1 U206 ( .A1(n2689), .A2(n2654), .ZN(n2667) );
  NOR3_X1 U207 ( .A1(n5710), .A2(n5707), .A3(n5720), .ZN(n5714) );
  NAND2_X1 U208 ( .A1(n2673), .A2(n2666), .ZN(n20267) );
  NAND2_X1 U209 ( .A1(n2673), .A2(n2666), .ZN(n20268) );
  NAND2_X1 U210 ( .A1(n5695), .A2(n5703), .ZN(n20082) );
  NAND2_X1 U211 ( .A1(n5695), .A2(n5703), .ZN(n20081) );
  NAND2_X1 U212 ( .A1(n2673), .A2(n2666), .ZN(n1861) );
  NAND2_X1 U213 ( .A1(n5699), .A2(n5700), .ZN(n20099) );
  NAND2_X1 U214 ( .A1(n5699), .A2(n5700), .ZN(n20098) );
  NOR3_X1 U215 ( .A1(n2675), .A2(n2653), .A3(n2690), .ZN(n2687) );
  NAND2_X1 U216 ( .A1(n5699), .A2(n5703), .ZN(n20048) );
  NAND2_X1 U217 ( .A1(n5699), .A2(n5703), .ZN(n20047) );
  NAND2_X1 U218 ( .A1(n5695), .A2(n5703), .ZN(n2713) );
  NAND2_X1 U219 ( .A1(n5699), .A2(n5700), .ZN(n2708) );
  NAND2_X1 U220 ( .A1(n5699), .A2(n5703), .ZN(n2717) );
  NAND2_X1 U221 ( .A1(n2674), .A2(n2673), .ZN(n20285) );
  NAND2_X1 U222 ( .A1(n2674), .A2(n2673), .ZN(n20286) );
  AND2_X1 U223 ( .A1(n2665), .A2(n2674), .ZN(n20294) );
  AND2_X1 U224 ( .A1(n2665), .A2(n2674), .ZN(n20295) );
  AND2_X1 U225 ( .A1(n2667), .A2(n2668), .ZN(n20313) );
  AND2_X1 U226 ( .A1(n2667), .A2(n2668), .ZN(n20314) );
  AND2_X1 U227 ( .A1(n5697), .A2(n5698), .ZN(n20101) );
  AND2_X1 U228 ( .A1(n5697), .A2(n5698), .ZN(n20100) );
  AND2_X1 U229 ( .A1(n2673), .A2(n2669), .ZN(n20296) );
  AND2_X1 U230 ( .A1(n2673), .A2(n2669), .ZN(n20297) );
  AND2_X1 U231 ( .A1(n5695), .A2(n5696), .ZN(n20103) );
  AND2_X1 U232 ( .A1(n5695), .A2(n5696), .ZN(n20102) );
  AND2_X1 U233 ( .A1(n2665), .A2(n2666), .ZN(n20315) );
  AND2_X1 U234 ( .A1(n2665), .A2(n2666), .ZN(n20316) );
  NAND2_X1 U235 ( .A1(n2674), .A2(n2673), .ZN(n1853) );
  AND2_X1 U236 ( .A1(n2665), .A2(n2674), .ZN(n1856) );
  AND2_X1 U237 ( .A1(n2667), .A2(n2668), .ZN(n1851) );
  AND2_X1 U238 ( .A1(n5697), .A2(n5698), .ZN(n2710) );
  AND2_X1 U239 ( .A1(n2673), .A2(n2669), .ZN(n1858) );
  AND2_X1 U240 ( .A1(n5695), .A2(n5696), .ZN(n2711) );
  AND2_X1 U241 ( .A1(n2665), .A2(n2666), .ZN(n1852) );
  AND2_X1 U242 ( .A1(n5695), .A2(n5698), .ZN(n2715) );
  AND2_X1 U243 ( .A1(n5695), .A2(n5698), .ZN(n20083) );
  NAND2_X1 U244 ( .A1(n5699), .A2(n5698), .ZN(n2712) );
  NOR2_X1 U245 ( .A1(n19781), .A2(n2696), .ZN(n2693) );
  NOR2_X1 U246 ( .A1(n20670), .A2(n1837), .ZN(n1834) );
  NAND2_X1 U247 ( .A1(n2665), .A2(n2669), .ZN(n1848) );
  NAND2_X1 U248 ( .A1(n2669), .A2(n2668), .ZN(n1865) );
  NAND2_X1 U249 ( .A1(n5703), .A2(n5706), .ZN(n2723) );
  NAND2_X1 U250 ( .A1(n5696), .A2(n5706), .ZN(n2724) );
  NAND2_X1 U251 ( .A1(n2665), .A2(n2667), .ZN(n20306) );
  NAND2_X1 U252 ( .A1(n2665), .A2(n2667), .ZN(n1849) );
  NAND2_X1 U253 ( .A1(n2676), .A2(n2666), .ZN(n1860) );
  NAND2_X1 U254 ( .A1(n2685), .A2(n2666), .ZN(n1878) );
  NAND2_X1 U255 ( .A1(n2685), .A2(n2669), .ZN(n1875) );
  NAND2_X1 U256 ( .A1(n2685), .A2(n2667), .ZN(n1892) );
  NAND2_X1 U257 ( .A1(n2685), .A2(n2674), .ZN(n1891) );
  NAND2_X1 U258 ( .A1(n2680), .A2(n2669), .ZN(n1866) );
  NAND2_X1 U259 ( .A1(n2687), .A2(n2669), .ZN(n1877) );
  NAND2_X1 U260 ( .A1(n2684), .A2(n2669), .ZN(n1885) );
  NAND2_X1 U261 ( .A1(n2687), .A2(n2666), .ZN(n1886) );
  NAND2_X1 U262 ( .A1(n5714), .A2(n5700), .ZN(n2734) );
  NAND2_X1 U263 ( .A1(n5717), .A2(n5698), .ZN(n2735) );
  NAND2_X1 U264 ( .A1(n5714), .A2(n5698), .ZN(n2732) );
  NAND2_X1 U265 ( .A1(n5717), .A2(n5700), .ZN(n2744) );
  NAND2_X1 U266 ( .A1(n5717), .A2(n5696), .ZN(n2749) );
  NAND2_X1 U267 ( .A1(n5714), .A2(n5696), .ZN(n2748) );
  NAND2_X1 U268 ( .A1(n2676), .A2(n2669), .ZN(n20287) );
  NAND2_X1 U269 ( .A1(n2676), .A2(n2669), .ZN(n1854) );
  NAND2_X1 U270 ( .A1(n5713), .A2(n5696), .ZN(n2743) );
  NAND2_X1 U271 ( .A1(n5713), .A2(n5698), .ZN(n2733) );
  NAND2_X1 U272 ( .A1(n2684), .A2(n2667), .ZN(n1876) );
  NAND2_X1 U273 ( .A1(n5701), .A2(n5696), .ZN(n20091) );
  NAND2_X1 U274 ( .A1(n5701), .A2(n5696), .ZN(n2707) );
  NAND2_X1 U275 ( .A1(n5700), .A2(n5706), .ZN(n2718) );
  AND2_X1 U276 ( .A1(n2673), .A2(n2667), .ZN(n1863) );
  AND2_X1 U277 ( .A1(n5699), .A2(n5696), .ZN(n2720) );
  AND2_X1 U278 ( .A1(n2666), .A2(n2668), .ZN(n1868) );
  AND2_X1 U279 ( .A1(n2666), .A2(n2680), .ZN(n1881) );
  AND2_X1 U280 ( .A1(n2667), .A2(n2676), .ZN(n1870) );
  AND2_X1 U281 ( .A1(n2667), .A2(n2680), .ZN(n1880) );
  AND2_X1 U282 ( .A1(n2684), .A2(n2666), .ZN(n1883) );
  AND2_X1 U283 ( .A1(n2674), .A2(n2676), .ZN(n1864) );
  AND2_X1 U284 ( .A1(n2674), .A2(n2680), .ZN(n1889) );
  AND2_X1 U285 ( .A1(n5717), .A2(n5703), .ZN(n2738) );
  AND2_X1 U286 ( .A1(n5713), .A2(n5703), .ZN(n2729) );
  AND2_X1 U287 ( .A1(n5697), .A2(n5703), .ZN(n2746) );
  AND2_X1 U288 ( .A1(n5714), .A2(n5703), .ZN(n2745) );
  AND2_X1 U289 ( .A1(n5697), .A2(n5696), .ZN(n2737) );
  AND2_X1 U290 ( .A1(n2684), .A2(n2674), .ZN(n1871) );
  AND2_X1 U291 ( .A1(n2687), .A2(n2674), .ZN(n1887) );
  AND2_X1 U292 ( .A1(n5701), .A2(n5698), .ZN(n2721) );
  AND2_X1 U293 ( .A1(n5713), .A2(n5700), .ZN(n2741) );
  AND2_X1 U294 ( .A1(n5701), .A2(n5700), .ZN(n2740) );
  AND2_X1 U295 ( .A1(n5698), .A2(n5706), .ZN(n2726) );
  AND2_X1 U296 ( .A1(n5700), .A2(n5695), .ZN(n20040) );
  AND2_X1 U297 ( .A1(n5700), .A2(n5695), .ZN(n2727) );
  INV_X1 U298 ( .A(n20532), .ZN(n1227) );
  INV_X1 U299 ( .A(n20534), .ZN(n1189) );
  AND2_X1 U300 ( .A1(n5697), .A2(n5700), .ZN(n20084) );
  AND2_X1 U301 ( .A1(n5697), .A2(n5700), .ZN(n2716) );
  INV_X1 U302 ( .A(n1439), .ZN(n20464) );
  INV_X1 U303 ( .A(n1371), .ZN(n20480) );
  INV_X1 U304 ( .A(n1657), .ZN(n20374) );
  INV_X1 U305 ( .A(n1446), .ZN(n20446) );
  INV_X1 U306 ( .A(n1297), .ZN(n20514) );
  INV_X1 U307 ( .A(n1263), .ZN(n20523) );
  BUF_X1 U308 ( .A(n20668), .Z(n20679) );
  INV_X1 U309 ( .A(n1335), .ZN(n20496) );
  BUF_X1 U310 ( .A(n1079), .Z(n20665) );
  BUF_X1 U311 ( .A(n20668), .Z(n20678) );
  BUF_X1 U312 ( .A(n20668), .Z(n20677) );
  BUF_X1 U313 ( .A(n20667), .Z(n20676) );
  BUF_X1 U314 ( .A(n20667), .Z(n20675) );
  BUF_X1 U315 ( .A(n20667), .Z(n20674) );
  BUF_X1 U316 ( .A(n20666), .Z(n20673) );
  BUF_X1 U317 ( .A(n20666), .Z(n20672) );
  BUF_X1 U318 ( .A(n20666), .Z(n20671) );
  INV_X1 U319 ( .A(n19889), .ZN(n2695) );
  BUF_X1 U320 ( .A(n1191), .Z(n19891) );
  BUF_X1 U321 ( .A(n1191), .Z(n19890) );
  BUF_X1 U322 ( .A(n1191), .Z(n19892) );
  NAND2_X1 U323 ( .A1(n1444), .A2(n1225), .ZN(n1554) );
  BUF_X1 U324 ( .A(n1187), .Z(n19894) );
  BUF_X1 U325 ( .A(n1187), .Z(n19893) );
  BUF_X1 U326 ( .A(n1187), .Z(n19895) );
  BUF_X1 U327 ( .A(n1079), .Z(n20664) );
  BUF_X1 U328 ( .A(n1079), .Z(n20663) );
  BUF_X1 U329 ( .A(n1079), .Z(n20662) );
  BUF_X1 U330 ( .A(n1079), .Z(n20661) );
  BUF_X1 U331 ( .A(n1079), .Z(n20660) );
  BUF_X1 U332 ( .A(n1079), .Z(n20659) );
  INV_X1 U333 ( .A(n1833), .ZN(n20320) );
  INV_X1 U334 ( .A(n1833), .ZN(n20321) );
  INV_X1 U335 ( .A(n1799), .ZN(n20329) );
  INV_X1 U336 ( .A(n1799), .ZN(n20330) );
  INV_X1 U337 ( .A(n1764), .ZN(n20338) );
  INV_X1 U338 ( .A(n1764), .ZN(n20339) );
  INV_X1 U339 ( .A(n1730), .ZN(n20347) );
  INV_X1 U340 ( .A(n1730), .ZN(n20348) );
  INV_X1 U341 ( .A(n1589), .ZN(n20392) );
  INV_X1 U342 ( .A(n1589), .ZN(n20393) );
  INV_X1 U343 ( .A(n1520), .ZN(n20410) );
  INV_X1 U344 ( .A(n1520), .ZN(n20411) );
  INV_X1 U345 ( .A(n1517), .ZN(n20419) );
  INV_X1 U346 ( .A(n1371), .ZN(n20481) );
  INV_X1 U347 ( .A(n1623), .ZN(n20383) );
  INV_X1 U348 ( .A(n1623), .ZN(n20384) );
  INV_X1 U349 ( .A(n1443), .ZN(n20455) );
  INV_X1 U350 ( .A(n1263), .ZN(n20524) );
  INV_X1 U351 ( .A(n1695), .ZN(n20356) );
  INV_X1 U352 ( .A(n1695), .ZN(n20357) );
  INV_X1 U353 ( .A(n1661), .ZN(n20365) );
  INV_X1 U354 ( .A(n1661), .ZN(n20366) );
  INV_X1 U355 ( .A(n1484), .ZN(n20428) );
  INV_X1 U356 ( .A(n1484), .ZN(n20429) );
  INV_X1 U357 ( .A(n1450), .ZN(n20437) );
  INV_X1 U358 ( .A(n1450), .ZN(n20438) );
  INV_X1 U359 ( .A(n1335), .ZN(n20497) );
  INV_X1 U360 ( .A(n1301), .ZN(n20505) );
  INV_X1 U361 ( .A(n1301), .ZN(n20506) );
  BUF_X1 U362 ( .A(n20489), .Z(n20490) );
  BUF_X1 U363 ( .A(n20489), .Z(n20491) );
  BUF_X1 U364 ( .A(n20489), .Z(n20492) );
  BUF_X1 U365 ( .A(n20473), .Z(n20474) );
  BUF_X1 U366 ( .A(n20473), .Z(n20475) );
  BUF_X1 U367 ( .A(n20473), .Z(n20476) );
  BUF_X1 U368 ( .A(n1368), .Z(n20493) );
  BUF_X1 U369 ( .A(n1368), .Z(n20494) );
  BUF_X1 U370 ( .A(n1405), .Z(n20477) );
  BUF_X1 U371 ( .A(n1405), .Z(n20478) );
  BUF_X1 U372 ( .A(n1368), .Z(n20495) );
  BUF_X1 U373 ( .A(n1405), .Z(n20479) );
  BUF_X1 U374 ( .A(n1148), .Z(n20549) );
  BUF_X1 U375 ( .A(n1148), .Z(n20548) );
  BUF_X1 U376 ( .A(n1148), .Z(n20547) );
  NAND2_X1 U377 ( .A1(n20686), .A2(n19881), .ZN(n18776) );
  NAND2_X1 U378 ( .A1(n20686), .A2(n19873), .ZN(n18773) );
  NAND2_X1 U379 ( .A1(n5683), .A2(n19876), .ZN(n3085) );
  NAND2_X1 U380 ( .A1(n5639), .A2(n19876), .ZN(n3097) );
  NAND2_X1 U381 ( .A1(n4950), .A2(n19876), .ZN(n3109) );
  NAND2_X1 U382 ( .A1(n4739), .A2(n19877), .ZN(n3133) );
  NAND2_X1 U383 ( .A1(n4695), .A2(n19878), .ZN(n3145) );
  NAND2_X1 U384 ( .A1(n4629), .A2(n19877), .ZN(n3163) );
  NAND2_X1 U385 ( .A1(n4607), .A2(n19878), .ZN(n3169) );
  NAND2_X1 U386 ( .A1(n4541), .A2(n19878), .ZN(n3187) );
  NAND2_X1 U387 ( .A1(n2927), .A2(n19876), .ZN(n3217) );
  NAND2_X1 U388 ( .A1(n2883), .A2(n19876), .ZN(n3229) );
  NAND2_X1 U389 ( .A1(n2861), .A2(n19877), .ZN(n3235) );
  NAND2_X1 U390 ( .A1(n2795), .A2(n19878), .ZN(n3253) );
  NAND2_X1 U391 ( .A1(n2773), .A2(n19878), .ZN(n3259) );
  NAND2_X1 U392 ( .A1(n5661), .A2(n19877), .ZN(n3091) );
  NAND2_X1 U393 ( .A1(n4915), .A2(n19878), .ZN(n3115) );
  NAND2_X1 U394 ( .A1(n4717), .A2(n19877), .ZN(n3139) );
  NAND2_X1 U395 ( .A1(n4651), .A2(n19876), .ZN(n3157) );
  NAND2_X1 U396 ( .A1(n2817), .A2(n19877), .ZN(n3247) );
  NAND2_X1 U397 ( .A1(n2644), .A2(n19868), .ZN(n3275) );
  NAND2_X1 U398 ( .A1(n2619), .A2(n19869), .ZN(n3280) );
  NAND2_X1 U399 ( .A1(n2594), .A2(n19868), .ZN(n3285) );
  NAND2_X1 U400 ( .A1(n2544), .A2(n19868), .ZN(n3295) );
  NAND2_X1 U401 ( .A1(n2519), .A2(n19870), .ZN(n3300) );
  NAND2_X1 U402 ( .A1(n2444), .A2(n19869), .ZN(n3315) );
  NAND2_X1 U403 ( .A1(n2419), .A2(n19869), .ZN(n3320) );
  NAND2_X1 U404 ( .A1(n2394), .A2(n19870), .ZN(n3325) );
  NAND2_X1 U405 ( .A1(n2344), .A2(n19868), .ZN(n3335) );
  NAND2_X1 U406 ( .A1(n2319), .A2(n19869), .ZN(n3340) );
  NAND2_X1 U407 ( .A1(n2294), .A2(n19870), .ZN(n3345) );
  NAND2_X1 U408 ( .A1(n2219), .A2(n19870), .ZN(n3360) );
  NAND2_X1 U409 ( .A1(n2094), .A2(n19868), .ZN(n3385) );
  NAND2_X1 U410 ( .A1(n2044), .A2(n19868), .ZN(n3395) );
  NAND2_X1 U411 ( .A1(n2019), .A2(n19869), .ZN(n3400) );
  NAND2_X1 U412 ( .A1(n1969), .A2(n19869), .ZN(n3410) );
  NAND2_X1 U413 ( .A1(n1944), .A2(n19870), .ZN(n3415) );
  NAND2_X1 U414 ( .A1(n1919), .A2(n19870), .ZN(n3420) );
  NAND2_X1 U415 ( .A1(n4879), .A2(n19879), .ZN(n3121) );
  NAND2_X1 U416 ( .A1(n4761), .A2(n19880), .ZN(n3127) );
  NAND2_X1 U417 ( .A1(n4585), .A2(n19879), .ZN(n3175) );
  NAND2_X1 U418 ( .A1(n4519), .A2(n19879), .ZN(n3193) );
  NAND2_X1 U419 ( .A1(n4497), .A2(n19880), .ZN(n3199) );
  NAND2_X1 U420 ( .A1(n4475), .A2(n19879), .ZN(n3205) );
  NAND2_X1 U421 ( .A1(n2839), .A2(n19880), .ZN(n3241) );
  NAND2_X1 U422 ( .A1(n2694), .A2(n19880), .ZN(n3271) );
  NAND2_X1 U423 ( .A1(n4563), .A2(n19880), .ZN(n3181) );
  NAND2_X1 U424 ( .A1(n2751), .A2(n19879), .ZN(n3265) );
  NAND2_X1 U425 ( .A1(n2494), .A2(n19871), .ZN(n3305) );
  NAND2_X1 U426 ( .A1(n2469), .A2(n19872), .ZN(n3310) );
  NAND2_X1 U427 ( .A1(n2269), .A2(n19871), .ZN(n3350) );
  NAND2_X1 U428 ( .A1(n2244), .A2(n19872), .ZN(n3355) );
  NAND2_X1 U429 ( .A1(n2194), .A2(n19871), .ZN(n3365) );
  NAND2_X1 U430 ( .A1(n2169), .A2(n19872), .ZN(n3370) );
  NAND2_X1 U431 ( .A1(n2144), .A2(n19871), .ZN(n3375) );
  NAND2_X1 U432 ( .A1(n1994), .A2(n19872), .ZN(n3405) );
  NAND2_X1 U433 ( .A1(n1894), .A2(n19871), .ZN(n3425) );
  NAND2_X1 U434 ( .A1(n1835), .A2(n19872), .ZN(n3430) );
  NAND2_X1 U435 ( .A1(n5321), .A2(n19881), .ZN(n3103) );
  NAND2_X1 U436 ( .A1(n4673), .A2(n19881), .ZN(n3151) );
  NAND2_X1 U437 ( .A1(n2949), .A2(n19881), .ZN(n3211) );
  NAND2_X1 U438 ( .A1(n2905), .A2(n19881), .ZN(n3223) );
  NAND2_X1 U439 ( .A1(n2569), .A2(n19873), .ZN(n3290) );
  NAND2_X1 U440 ( .A1(n2369), .A2(n19873), .ZN(n3330) );
  NAND2_X1 U441 ( .A1(n2119), .A2(n19873), .ZN(n3380) );
  NAND2_X1 U442 ( .A1(n2069), .A2(n19873), .ZN(n3390) );
  INV_X2 U443 ( .A(n5684), .ZN(n2696) );
  INV_X2 U444 ( .A(n2645), .ZN(n1837) );
  NOR3_X1 U445 ( .A1(n5710), .A2(ADD_RD1[0]), .A3(n5720), .ZN(n5697) );
  NOR3_X1 U446 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n2653), .ZN(n2676) );
  NOR3_X1 U447 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n2690), .ZN(n2685) );
  NOR3_X1 U448 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n5710), .ZN(n5706) );
  NOR3_X1 U449 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(n2668)
         );
  NOR3_X1 U450 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n5720), .ZN(n5717) );
  NOR3_X1 U451 ( .A1(n5707), .A2(ADD_RD1[3]), .A3(n5720), .ZN(n5713) );
  NOR3_X1 U452 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(n5701)
         );
  NOR3_X1 U453 ( .A1(n2653), .A2(ADD_RD2[3]), .A3(n2690), .ZN(n2684) );
  NAND2_X1 U454 ( .A1(n1225), .A2(n1145), .ZN(n20532) );
  NAND2_X1 U455 ( .A1(n1188), .A2(n1145), .ZN(n20534) );
  NOR3_X1 U456 ( .A1(n2675), .A2(ADD_RD2[0]), .A3(n2690), .ZN(n2680) );
  AND2_X1 U457 ( .A1(ADD_RD1[2]), .A2(ADD_RD1[1]), .ZN(n5700) );
  AND2_X1 U458 ( .A1(ADD_RD1[2]), .A2(n5718), .ZN(n5698) );
  OAI22_X1 U459 ( .A1(n19235), .A2(n19946), .B1(n18883), .B2(n19953), .ZN(
        n5719) );
  OAI22_X1 U460 ( .A1(n18851), .A2(n19914), .B1(n19107), .B2(n19922), .ZN(
        n5721) );
  OAI22_X1 U461 ( .A1(n19237), .A2(n19951), .B1(n18885), .B2(n19959), .ZN(
        n5659) );
  OAI22_X1 U462 ( .A1(n18853), .A2(n19917), .B1(n19109), .B2(n19927), .ZN(
        n5660) );
  OAI22_X1 U463 ( .A1(n19238), .A2(n19951), .B1(n18886), .B2(n19956), .ZN(
        n5637) );
  OAI22_X1 U464 ( .A1(n18854), .A2(n19917), .B1(n19110), .B2(n19926), .ZN(
        n5638) );
  OAI22_X1 U465 ( .A1(n19239), .A2(n19951), .B1(n18887), .B2(n19958), .ZN(
        n5319) );
  OAI22_X1 U466 ( .A1(n18855), .A2(n19917), .B1(n19111), .B2(n19927), .ZN(
        n5320) );
  OAI22_X1 U467 ( .A1(n19241), .A2(n19947), .B1(n18889), .B2(n19954), .ZN(
        n4913) );
  OAI22_X1 U468 ( .A1(n18857), .A2(n19915), .B1(n19113), .B2(n19923), .ZN(
        n4914) );
  OAI22_X1 U469 ( .A1(n19242), .A2(n19948), .B1(n18890), .B2(n19955), .ZN(
        n4877) );
  OAI22_X1 U470 ( .A1(n18858), .A2(n19916), .B1(n19114), .B2(n19924), .ZN(
        n4878) );
  OAI22_X1 U471 ( .A1(n19243), .A2(n19950), .B1(n18891), .B2(n19956), .ZN(
        n4759) );
  OAI22_X1 U472 ( .A1(n18859), .A2(n19918), .B1(n19115), .B2(n19925), .ZN(
        n4760) );
  OAI22_X1 U473 ( .A1(n19245), .A2(n19949), .B1(n18893), .B2(n19956), .ZN(
        n4715) );
  OAI22_X1 U474 ( .A1(n18861), .A2(n19917), .B1(n19117), .B2(n19925), .ZN(
        n4716) );
  OAI22_X1 U475 ( .A1(n19246), .A2(n19950), .B1(n18894), .B2(n19957), .ZN(
        n4693) );
  OAI22_X1 U476 ( .A1(n18862), .A2(n19918), .B1(n19118), .B2(n19926), .ZN(
        n4694) );
  OAI22_X1 U477 ( .A1(n19248), .A2(n19946), .B1(n18896), .B2(n19953), .ZN(
        n4649) );
  OAI22_X1 U478 ( .A1(n18864), .A2(n19915), .B1(n19120), .B2(n19923), .ZN(
        n4650) );
  OAI22_X1 U479 ( .A1(n19249), .A2(n19947), .B1(n18897), .B2(n19954), .ZN(
        n4627) );
  OAI22_X1 U480 ( .A1(n18865), .A2(n19915), .B1(n19121), .B2(n19923), .ZN(
        n4628) );
  OAI22_X1 U481 ( .A1(n19250), .A2(n19948), .B1(n18898), .B2(n19955), .ZN(
        n4605) );
  OAI22_X1 U482 ( .A1(n18866), .A2(n19916), .B1(n19122), .B2(n19924), .ZN(
        n4606) );
  OAI22_X1 U483 ( .A1(n19252), .A2(n19946), .B1(n18900), .B2(n19955), .ZN(
        n4561) );
  OAI22_X1 U484 ( .A1(n18868), .A2(n19915), .B1(n19124), .B2(n19922), .ZN(
        n4562) );
  OAI22_X1 U485 ( .A1(n19253), .A2(n19949), .B1(n18901), .B2(n19956), .ZN(
        n4539) );
  OAI22_X1 U486 ( .A1(n18869), .A2(n19917), .B1(n19125), .B2(n19925), .ZN(
        n4540) );
  OAI22_X1 U487 ( .A1(n19254), .A2(n19950), .B1(n18902), .B2(n19957), .ZN(
        n4517) );
  OAI22_X1 U488 ( .A1(n18870), .A2(n19918), .B1(n19126), .B2(n19926), .ZN(
        n4518) );
  OAI22_X1 U489 ( .A1(n19255), .A2(n19946), .B1(n18903), .B2(n19954), .ZN(
        n2815) );
  OAI22_X1 U490 ( .A1(n18871), .A2(n19914), .B1(n19135), .B2(n19924), .ZN(
        n2816) );
  OAI22_X1 U491 ( .A1(n19256), .A2(n19948), .B1(n18904), .B2(n19953), .ZN(
        n2793) );
  OAI22_X1 U492 ( .A1(n18872), .A2(n19916), .B1(n19136), .B2(n19922), .ZN(
        n2794) );
  OAI22_X1 U493 ( .A1(n19258), .A2(n19950), .B1(n18906), .B2(n19958), .ZN(
        n2742) );
  OAI22_X1 U494 ( .A1(n18874), .A2(n19918), .B1(n19138), .B2(n19925), .ZN(
        n2747) );
  OAI22_X1 U495 ( .A1(n19236), .A2(n19947), .B1(n18884), .B2(n19953), .ZN(
        n5681) );
  OAI22_X1 U496 ( .A1(n18852), .A2(n19914), .B1(n19108), .B2(n19922), .ZN(
        n5682) );
  OAI22_X1 U497 ( .A1(n19240), .A2(n19948), .B1(n18888), .B2(n19955), .ZN(
        n4948) );
  OAI22_X1 U498 ( .A1(n18856), .A2(n19914), .B1(n19112), .B2(n19924), .ZN(
        n4949) );
  OAI22_X1 U499 ( .A1(n19244), .A2(n19947), .B1(n18892), .B2(n19954), .ZN(
        n4737) );
  OAI22_X1 U500 ( .A1(n18860), .A2(n19916), .B1(n19116), .B2(n19923), .ZN(
        n4738) );
  OAI22_X1 U501 ( .A1(n19247), .A2(n19949), .B1(n18895), .B2(n19956), .ZN(
        n4671) );
  OAI22_X1 U502 ( .A1(n18863), .A2(n19918), .B1(n19119), .B2(n19925), .ZN(
        n4672) );
  OAI22_X1 U503 ( .A1(n19251), .A2(n19950), .B1(n18899), .B2(n19959), .ZN(
        n4583) );
  OAI22_X1 U504 ( .A1(n18867), .A2(n19919), .B1(n19123), .B2(n19926), .ZN(
        n4584) );
  OAI22_X1 U505 ( .A1(n19257), .A2(n19949), .B1(n18905), .B2(n19957), .ZN(
        n2771) );
  OAI22_X1 U506 ( .A1(n18873), .A2(n19919), .B1(n19137), .B2(n19926), .ZN(
        n2772) );
  OAI22_X1 U507 ( .A1(n19043), .A2(n20162), .B1(n18851), .B2(n20164), .ZN(
        n2688) );
  OAI22_X1 U508 ( .A1(n19044), .A2(n20161), .B1(n18852), .B2(n20169), .ZN(
        n2640) );
  OAI22_X1 U509 ( .A1(n19045), .A2(n20161), .B1(n18853), .B2(n20169), .ZN(
        n2615) );
  OAI22_X1 U510 ( .A1(n19046), .A2(n20161), .B1(n18854), .B2(n20164), .ZN(
        n2590) );
  OAI22_X1 U511 ( .A1(n19047), .A2(n20156), .B1(n18855), .B2(n20165), .ZN(
        n2565) );
  OAI22_X1 U512 ( .A1(n19048), .A2(n20158), .B1(n18856), .B2(n20166), .ZN(
        n2540) );
  OAI22_X1 U513 ( .A1(n19049), .A2(n20157), .B1(n18857), .B2(n20165), .ZN(
        n2515) );
  OAI22_X1 U514 ( .A1(n19050), .A2(n20157), .B1(n18858), .B2(n20167), .ZN(
        n2490) );
  OAI22_X1 U515 ( .A1(n19051), .A2(n20156), .B1(n18859), .B2(n20167), .ZN(
        n2465) );
  OAI22_X1 U516 ( .A1(n19052), .A2(n20158), .B1(n18860), .B2(n20165), .ZN(
        n2440) );
  OAI22_X1 U517 ( .A1(n19053), .A2(n20160), .B1(n18861), .B2(n20170), .ZN(
        n2415) );
  OAI22_X1 U518 ( .A1(n19054), .A2(n20159), .B1(n18862), .B2(n20168), .ZN(
        n2390) );
  OAI22_X1 U519 ( .A1(n19055), .A2(n20156), .B1(n18863), .B2(n20165), .ZN(
        n2365) );
  OAI22_X1 U520 ( .A1(n19056), .A2(n20157), .B1(n18864), .B2(n20166), .ZN(
        n2340) );
  OAI22_X1 U521 ( .A1(n19057), .A2(n20157), .B1(n18865), .B2(n20166), .ZN(
        n2315) );
  OAI22_X1 U522 ( .A1(n19058), .A2(n20156), .B1(n18866), .B2(n20166), .ZN(
        n2290) );
  OAI22_X1 U523 ( .A1(n19059), .A2(n20157), .B1(n18867), .B2(n20167), .ZN(
        n2265) );
  OAI22_X1 U524 ( .A1(n19060), .A2(n20158), .B1(n18868), .B2(n20167), .ZN(
        n2240) );
  OAI22_X1 U525 ( .A1(n19061), .A2(n20162), .B1(n18869), .B2(n20169), .ZN(
        n2215) );
  OAI22_X1 U526 ( .A1(n19062), .A2(n20159), .B1(n18870), .B2(n20168), .ZN(
        n2190) );
  OAI22_X1 U527 ( .A1(n19063), .A2(n20158), .B1(n18875), .B2(n20164), .ZN(
        n2165) );
  OAI22_X1 U528 ( .A1(n19064), .A2(n20160), .B1(n18876), .B2(n20169), .ZN(
        n2140) );
  OAI22_X1 U529 ( .A1(n19065), .A2(n20161), .B1(n18877), .B2(n20170), .ZN(
        n2115) );
  OAI22_X1 U530 ( .A1(n19066), .A2(n20160), .B1(n18881), .B2(n20169), .ZN(
        n2090) );
  OAI22_X1 U531 ( .A1(n19067), .A2(n20161), .B1(n18878), .B2(n20170), .ZN(
        n2065) );
  OAI22_X1 U532 ( .A1(n19068), .A2(n20162), .B1(n18879), .B2(n20168), .ZN(
        n2040) );
  OAI22_X1 U533 ( .A1(n19069), .A2(n20162), .B1(n18880), .B2(n20170), .ZN(
        n2015) );
  OAI22_X1 U534 ( .A1(n19070), .A2(n20156), .B1(n18882), .B2(n20164), .ZN(
        n1990) );
  OAI22_X1 U535 ( .A1(n19071), .A2(n20159), .B1(n18871), .B2(n20164), .ZN(
        n1965) );
  OAI22_X1 U536 ( .A1(n19072), .A2(n20160), .B1(n18872), .B2(n20164), .ZN(
        n1940) );
  OAI22_X1 U537 ( .A1(n19073), .A2(n20162), .B1(n18873), .B2(n20170), .ZN(
        n1915) );
  OAI22_X1 U538 ( .A1(n19074), .A2(n20159), .B1(n18874), .B2(n20168), .ZN(
        n1884) );
  OAI22_X1 U539 ( .A1(n18915), .A2(n20004), .B1(n19043), .B2(n20015), .ZN(
        n5712) );
  OAI22_X1 U540 ( .A1(n18917), .A2(n20007), .B1(n19045), .B2(n20012), .ZN(
        n5656) );
  OAI22_X1 U541 ( .A1(n18918), .A2(n20005), .B1(n19046), .B2(n20013), .ZN(
        n5634) );
  OAI22_X1 U542 ( .A1(n18919), .A2(n20002), .B1(n19047), .B2(n20010), .ZN(
        n5316) );
  OAI22_X1 U543 ( .A1(n18921), .A2(n20003), .B1(n19049), .B2(n20009), .ZN(
        n4910) );
  OAI22_X1 U544 ( .A1(n18922), .A2(n20004), .B1(n19050), .B2(n20009), .ZN(
        n4778) );
  OAI22_X1 U545 ( .A1(n18923), .A2(n20001), .B1(n19051), .B2(n20012), .ZN(
        n4756) );
  OAI22_X1 U546 ( .A1(n18925), .A2(n20005), .B1(n19053), .B2(n20010), .ZN(
        n4712) );
  OAI22_X1 U547 ( .A1(n18926), .A2(n20006), .B1(n19054), .B2(n20011), .ZN(
        n4690) );
  OAI22_X1 U548 ( .A1(n18928), .A2(n20002), .B1(n19056), .B2(n20010), .ZN(
        n4646) );
  OAI22_X1 U549 ( .A1(n18929), .A2(n20003), .B1(n19057), .B2(n20009), .ZN(
        n4624) );
  OAI22_X1 U550 ( .A1(n18930), .A2(n20004), .B1(n19058), .B2(n20009), .ZN(
        n4602) );
  OAI22_X1 U551 ( .A1(n18932), .A2(n20003), .B1(n19060), .B2(n20010), .ZN(
        n4558) );
  OAI22_X1 U552 ( .A1(n18933), .A2(n20005), .B1(n19061), .B2(n20010), .ZN(
        n4536) );
  OAI22_X1 U553 ( .A1(n18934), .A2(n20006), .B1(n19062), .B2(n20011), .ZN(
        n4514) );
  OAI22_X1 U554 ( .A1(n18935), .A2(n20006), .B1(n19063), .B2(n20012), .ZN(
        n4492) );
  OAI22_X1 U555 ( .A1(n18936), .A2(n20007), .B1(n19064), .B2(n20013), .ZN(
        n4470) );
  OAI22_X1 U556 ( .A1(n18937), .A2(n20007), .B1(n19065), .B2(n20013), .ZN(
        n2944) );
  OAI22_X1 U557 ( .A1(n18939), .A2(n20005), .B1(n19067), .B2(n20014), .ZN(
        n2900) );
  OAI22_X1 U558 ( .A1(n18940), .A2(n20002), .B1(n19068), .B2(n20014), .ZN(
        n2878) );
  OAI22_X1 U559 ( .A1(n18941), .A2(n20007), .B1(n19069), .B2(n20015), .ZN(
        n2856) );
  OAI22_X1 U560 ( .A1(n18943), .A2(n20003), .B1(n19071), .B2(n20014), .ZN(
        n2812) );
  OAI22_X1 U561 ( .A1(n18944), .A2(n20001), .B1(n19072), .B2(n20015), .ZN(
        n2790) );
  OAI22_X1 U562 ( .A1(n18946), .A2(n20006), .B1(n19074), .B2(n20011), .ZN(
        n2731) );
  OAI22_X1 U563 ( .A1(n18916), .A2(n20001), .B1(n19044), .B2(n20014), .ZN(
        n5678) );
  OAI22_X1 U564 ( .A1(n18920), .A2(n20002), .B1(n19048), .B2(n20012), .ZN(
        n4945) );
  OAI22_X1 U565 ( .A1(n18924), .A2(n20004), .B1(n19052), .B2(n20010), .ZN(
        n4734) );
  OAI22_X1 U566 ( .A1(n18927), .A2(n20002), .B1(n19055), .B2(n20011), .ZN(
        n4668) );
  OAI22_X1 U567 ( .A1(n18931), .A2(n20001), .B1(n19059), .B2(n20013), .ZN(
        n4580) );
  OAI22_X1 U568 ( .A1(n18938), .A2(n20005), .B1(n19066), .B2(n20015), .ZN(
        n2922) );
  OAI22_X1 U569 ( .A1(n18942), .A2(n20007), .B1(n19070), .B2(n20012), .ZN(
        n2834) );
  OAI22_X1 U570 ( .A1(n18945), .A2(n20005), .B1(n19073), .B2(n20013), .ZN(
        n2768) );
  BUF_X1 U571 ( .A(n1143), .Z(n20561) );
  BUF_X1 U572 ( .A(n1141), .Z(n20564) );
  BUF_X1 U573 ( .A(n1139), .Z(n20567) );
  BUF_X1 U574 ( .A(n1137), .Z(n20570) );
  BUF_X1 U575 ( .A(n1135), .Z(n20573) );
  BUF_X1 U576 ( .A(n1133), .Z(n20576) );
  BUF_X1 U577 ( .A(n1131), .Z(n20579) );
  BUF_X1 U578 ( .A(n1129), .Z(n20582) );
  BUF_X1 U579 ( .A(n1127), .Z(n20585) );
  BUF_X1 U580 ( .A(n1125), .Z(n20588) );
  BUF_X1 U581 ( .A(n1123), .Z(n20591) );
  BUF_X1 U582 ( .A(n1121), .Z(n20594) );
  BUF_X1 U583 ( .A(n1119), .Z(n20597) );
  BUF_X1 U584 ( .A(n1117), .Z(n20600) );
  BUF_X1 U585 ( .A(n1115), .Z(n20603) );
  BUF_X1 U586 ( .A(n1113), .Z(n20606) );
  BUF_X1 U587 ( .A(n1111), .Z(n20609) );
  BUF_X1 U588 ( .A(n1109), .Z(n20612) );
  BUF_X1 U589 ( .A(n1107), .Z(n20615) );
  BUF_X1 U590 ( .A(n1105), .Z(n20618) );
  BUF_X1 U591 ( .A(n1103), .Z(n20621) );
  BUF_X1 U592 ( .A(n1101), .Z(n20624) );
  BUF_X1 U593 ( .A(n1099), .Z(n20627) );
  BUF_X1 U594 ( .A(n1097), .Z(n20630) );
  BUF_X1 U595 ( .A(n1095), .Z(n20633) );
  BUF_X1 U596 ( .A(n1093), .Z(n20636) );
  BUF_X1 U597 ( .A(n1091), .Z(n20639) );
  BUF_X1 U598 ( .A(n1089), .Z(n20642) );
  BUF_X1 U599 ( .A(n1087), .Z(n20645) );
  BUF_X1 U600 ( .A(n1085), .Z(n20648) );
  BUF_X1 U601 ( .A(n1083), .Z(n20651) );
  BUF_X1 U602 ( .A(n1080), .Z(n20654) );
  BUF_X1 U603 ( .A(n1143), .Z(n20562) );
  BUF_X1 U604 ( .A(n1141), .Z(n20565) );
  BUF_X1 U605 ( .A(n1139), .Z(n20568) );
  BUF_X1 U606 ( .A(n1137), .Z(n20571) );
  BUF_X1 U607 ( .A(n1135), .Z(n20574) );
  BUF_X1 U608 ( .A(n1133), .Z(n20577) );
  BUF_X1 U609 ( .A(n1131), .Z(n20580) );
  BUF_X1 U610 ( .A(n1129), .Z(n20583) );
  BUF_X1 U611 ( .A(n1127), .Z(n20586) );
  BUF_X1 U612 ( .A(n1125), .Z(n20589) );
  BUF_X1 U613 ( .A(n1123), .Z(n20592) );
  BUF_X1 U614 ( .A(n1121), .Z(n20595) );
  BUF_X1 U615 ( .A(n1119), .Z(n20598) );
  BUF_X1 U616 ( .A(n1117), .Z(n20601) );
  BUF_X1 U617 ( .A(n1115), .Z(n20604) );
  BUF_X1 U618 ( .A(n1113), .Z(n20607) );
  BUF_X1 U619 ( .A(n1111), .Z(n20610) );
  BUF_X1 U620 ( .A(n1109), .Z(n20613) );
  BUF_X1 U621 ( .A(n1107), .Z(n20616) );
  BUF_X1 U622 ( .A(n1105), .Z(n20619) );
  BUF_X1 U623 ( .A(n1103), .Z(n20622) );
  BUF_X1 U624 ( .A(n1101), .Z(n20625) );
  BUF_X1 U625 ( .A(n1099), .Z(n20628) );
  BUF_X1 U626 ( .A(n1097), .Z(n20631) );
  BUF_X1 U627 ( .A(n1095), .Z(n20634) );
  BUF_X1 U628 ( .A(n1093), .Z(n20637) );
  BUF_X1 U629 ( .A(n1091), .Z(n20640) );
  BUF_X1 U630 ( .A(n1089), .Z(n20643) );
  BUF_X1 U631 ( .A(n1087), .Z(n20646) );
  BUF_X1 U632 ( .A(n1085), .Z(n20649) );
  BUF_X1 U633 ( .A(n1083), .Z(n20652) );
  BUF_X1 U634 ( .A(n1080), .Z(n20655) );
  OAI22_X1 U635 ( .A1(n20563), .A2(n20533), .B1(n19854), .B2(n19363), .ZN(
        n4171) );
  OAI22_X1 U636 ( .A1(n20566), .A2(n1226), .B1(n19854), .B2(n19379), .ZN(n4172) );
  OAI22_X1 U637 ( .A1(n20569), .A2(n20532), .B1(n19854), .B2(n19385), .ZN(
        n4173) );
  OAI22_X1 U638 ( .A1(n20572), .A2(n20533), .B1(n19854), .B2(n19364), .ZN(
        n4174) );
  OAI22_X1 U639 ( .A1(n20575), .A2(n1226), .B1(n19854), .B2(n19365), .ZN(n4175) );
  OAI22_X1 U640 ( .A1(n20578), .A2(n20532), .B1(n19854), .B2(n19393), .ZN(
        n4176) );
  OAI22_X1 U641 ( .A1(n20581), .A2(n20533), .B1(n19854), .B2(n19366), .ZN(
        n4177) );
  OAI22_X1 U642 ( .A1(n20584), .A2(n1226), .B1(n19854), .B2(n19367), .ZN(n4178) );
  OAI22_X1 U643 ( .A1(n20587), .A2(n20532), .B1(n19854), .B2(n19386), .ZN(
        n4179) );
  OAI22_X1 U644 ( .A1(n20590), .A2(n20533), .B1(n19854), .B2(n19380), .ZN(
        n4180) );
  OAI22_X1 U645 ( .A1(n20593), .A2(n1226), .B1(n19854), .B2(n19368), .ZN(n4181) );
  OAI22_X1 U646 ( .A1(n20596), .A2(n20532), .B1(n19854), .B2(n19387), .ZN(
        n4182) );
  OAI22_X1 U647 ( .A1(n20599), .A2(n20533), .B1(n19855), .B2(n19381), .ZN(
        n4183) );
  OAI22_X1 U648 ( .A1(n20602), .A2(n1226), .B1(n19855), .B2(n19369), .ZN(n4184) );
  OAI22_X1 U649 ( .A1(n20605), .A2(n20532), .B1(n19855), .B2(n19388), .ZN(
        n4185) );
  OAI22_X1 U650 ( .A1(n20608), .A2(n20533), .B1(n19855), .B2(n19370), .ZN(
        n4186) );
  OAI22_X1 U651 ( .A1(n20611), .A2(n1226), .B1(n19855), .B2(n19382), .ZN(n4187) );
  OAI22_X1 U652 ( .A1(n20614), .A2(n20532), .B1(n19855), .B2(n19389), .ZN(
        n4188) );
  OAI22_X1 U653 ( .A1(n20617), .A2(n20533), .B1(n19855), .B2(n19371), .ZN(
        n4189) );
  OAI22_X1 U654 ( .A1(n20620), .A2(n1226), .B1(n19855), .B2(n19372), .ZN(n4190) );
  OAI22_X1 U655 ( .A1(n20623), .A2(n20532), .B1(n19855), .B2(n19390), .ZN(
        n4191) );
  OAI22_X1 U656 ( .A1(n20626), .A2(n20533), .B1(n19855), .B2(n19373), .ZN(
        n4192) );
  OAI22_X1 U657 ( .A1(n20629), .A2(n1226), .B1(n19855), .B2(n19374), .ZN(n4193) );
  OAI22_X1 U658 ( .A1(n20632), .A2(n20532), .B1(n19855), .B2(n19394), .ZN(
        n4194) );
  NAND2_X1 U659 ( .A1(n1298), .A2(n1225), .ZN(n1439) );
  NAND2_X1 U660 ( .A1(n1298), .A2(n1188), .ZN(n1371) );
  OAI22_X1 U661 ( .A1(n20660), .A2(n20633), .B1(n20657), .B2(n19023), .ZN(
        n4387) );
  OAI22_X1 U662 ( .A1(n20660), .A2(n20636), .B1(n20658), .B2(n19024), .ZN(
        n4388) );
  OAI22_X1 U663 ( .A1(n20660), .A2(n20639), .B1(n20657), .B2(n19039), .ZN(
        n4389) );
  OAI22_X1 U664 ( .A1(n20659), .A2(n20642), .B1(n20658), .B2(n19031), .ZN(
        n4390) );
  OAI22_X1 U665 ( .A1(n20659), .A2(n20645), .B1(n20657), .B2(n19025), .ZN(
        n4391) );
  OAI22_X1 U666 ( .A1(n20659), .A2(n20648), .B1(n20658), .B2(n19040), .ZN(
        n4392) );
  OAI22_X1 U667 ( .A1(n20659), .A2(n20651), .B1(n20657), .B2(n19032), .ZN(
        n4393) );
  OAI22_X1 U668 ( .A1(n20659), .A2(n20654), .B1(n20658), .B2(n19026), .ZN(
        n4394) );
  OAI22_X1 U669 ( .A1(n20635), .A2(n20533), .B1(n19856), .B2(n19375), .ZN(
        n4195) );
  OAI22_X1 U670 ( .A1(n20638), .A2(n1226), .B1(n19856), .B2(n19376), .ZN(n4196) );
  OAI22_X1 U671 ( .A1(n20641), .A2(n20532), .B1(n19856), .B2(n19391), .ZN(
        n4197) );
  OAI22_X1 U672 ( .A1(n20644), .A2(n20533), .B1(n19856), .B2(n19383), .ZN(
        n4198) );
  OAI22_X1 U673 ( .A1(n20647), .A2(n1226), .B1(n19856), .B2(n19377), .ZN(n4199) );
  OAI22_X1 U674 ( .A1(n20650), .A2(n20532), .B1(n19856), .B2(n19392), .ZN(
        n4200) );
  OAI22_X1 U675 ( .A1(n20653), .A2(n20533), .B1(n19856), .B2(n19384), .ZN(
        n4201) );
  OAI22_X1 U676 ( .A1(n20656), .A2(n1226), .B1(n19856), .B2(n19378), .ZN(n4202) );
  OAI22_X1 U677 ( .A1(n20665), .A2(n20561), .B1(n20657), .B2(n19011), .ZN(
        n4363) );
  OAI22_X1 U678 ( .A1(n20665), .A2(n20564), .B1(n20657), .B2(n19027), .ZN(
        n4364) );
  OAI22_X1 U679 ( .A1(n20664), .A2(n20567), .B1(n20657), .B2(n19033), .ZN(
        n4365) );
  OAI22_X1 U680 ( .A1(n20664), .A2(n20570), .B1(n20657), .B2(n19012), .ZN(
        n4366) );
  OAI22_X1 U681 ( .A1(n20664), .A2(n20573), .B1(n20657), .B2(n19013), .ZN(
        n4367) );
  OAI22_X1 U682 ( .A1(n20664), .A2(n20576), .B1(n20657), .B2(n19041), .ZN(
        n4368) );
  OAI22_X1 U683 ( .A1(n20664), .A2(n20579), .B1(n20657), .B2(n19014), .ZN(
        n4369) );
  OAI22_X1 U684 ( .A1(n20663), .A2(n20582), .B1(n20657), .B2(n19015), .ZN(
        n4370) );
  OAI22_X1 U685 ( .A1(n20663), .A2(n20585), .B1(n20657), .B2(n19034), .ZN(
        n4371) );
  OAI22_X1 U686 ( .A1(n20663), .A2(n20588), .B1(n20657), .B2(n19028), .ZN(
        n4372) );
  OAI22_X1 U687 ( .A1(n20663), .A2(n20591), .B1(n20657), .B2(n19016), .ZN(
        n4373) );
  OAI22_X1 U688 ( .A1(n20663), .A2(n20594), .B1(n20657), .B2(n19035), .ZN(
        n4374) );
  OAI22_X1 U689 ( .A1(n20662), .A2(n20597), .B1(n20658), .B2(n19029), .ZN(
        n4375) );
  OAI22_X1 U690 ( .A1(n20662), .A2(n20600), .B1(n20658), .B2(n19017), .ZN(
        n4376) );
  OAI22_X1 U691 ( .A1(n20662), .A2(n20603), .B1(n20658), .B2(n19036), .ZN(
        n4377) );
  OAI22_X1 U692 ( .A1(n20662), .A2(n20606), .B1(n20658), .B2(n19018), .ZN(
        n4378) );
  OAI22_X1 U693 ( .A1(n20662), .A2(n20609), .B1(n20658), .B2(n19030), .ZN(
        n4379) );
  OAI22_X1 U694 ( .A1(n20661), .A2(n20612), .B1(n20658), .B2(n19037), .ZN(
        n4380) );
  OAI22_X1 U695 ( .A1(n20661), .A2(n20615), .B1(n20658), .B2(n19019), .ZN(
        n4381) );
  OAI22_X1 U696 ( .A1(n20661), .A2(n20618), .B1(n20658), .B2(n19020), .ZN(
        n4382) );
  OAI22_X1 U697 ( .A1(n20661), .A2(n20621), .B1(n20658), .B2(n19038), .ZN(
        n4383) );
  OAI22_X1 U698 ( .A1(n20661), .A2(n20624), .B1(n20658), .B2(n19021), .ZN(
        n4384) );
  OAI22_X1 U699 ( .A1(n20660), .A2(n20627), .B1(n20658), .B2(n19022), .ZN(
        n4385) );
  OAI22_X1 U700 ( .A1(n20660), .A2(n20630), .B1(n20658), .B2(n19042), .ZN(
        n4386) );
  OAI22_X1 U701 ( .A1(n19788), .A2(n18915), .B1(n20563), .B2(n20341), .ZN(
        n3467) );
  OAI22_X1 U702 ( .A1(n19788), .A2(n18916), .B1(n20566), .B2(n20340), .ZN(
        n3468) );
  OAI22_X1 U703 ( .A1(n19788), .A2(n18917), .B1(n20569), .B2(n20341), .ZN(
        n3469) );
  OAI22_X1 U704 ( .A1(n19788), .A2(n18918), .B1(n20572), .B2(n20343), .ZN(
        n3470) );
  OAI22_X1 U705 ( .A1(n19788), .A2(n18919), .B1(n20575), .B2(n20341), .ZN(
        n3471) );
  OAI22_X1 U706 ( .A1(n19788), .A2(n18920), .B1(n20578), .B2(n20346), .ZN(
        n3472) );
  OAI22_X1 U707 ( .A1(n19788), .A2(n18921), .B1(n20581), .B2(n20342), .ZN(
        n3473) );
  OAI22_X1 U708 ( .A1(n19788), .A2(n18922), .B1(n20584), .B2(n20343), .ZN(
        n3474) );
  OAI22_X1 U709 ( .A1(n19788), .A2(n18923), .B1(n20587), .B2(n20343), .ZN(
        n3475) );
  OAI22_X1 U710 ( .A1(n19788), .A2(n18924), .B1(n20590), .B2(n20345), .ZN(
        n3476) );
  OAI22_X1 U711 ( .A1(n19788), .A2(n18925), .B1(n20593), .B2(n20345), .ZN(
        n3477) );
  OAI22_X1 U712 ( .A1(n19788), .A2(n18926), .B1(n20596), .B2(n20344), .ZN(
        n3478) );
  OAI22_X1 U713 ( .A1(n19789), .A2(n18927), .B1(n20599), .B2(n20342), .ZN(
        n3479) );
  OAI22_X1 U714 ( .A1(n19789), .A2(n18928), .B1(n20602), .B2(n20343), .ZN(
        n3480) );
  OAI22_X1 U715 ( .A1(n19789), .A2(n18929), .B1(n20605), .B2(n20342), .ZN(
        n3481) );
  OAI22_X1 U716 ( .A1(n19789), .A2(n18930), .B1(n20608), .B2(n20344), .ZN(
        n3482) );
  OAI22_X1 U717 ( .A1(n19789), .A2(n18931), .B1(n20611), .B2(n20344), .ZN(
        n3483) );
  OAI22_X1 U718 ( .A1(n19789), .A2(n18932), .B1(n20614), .B2(n20344), .ZN(
        n3484) );
  OAI22_X1 U719 ( .A1(n19789), .A2(n18933), .B1(n20617), .B2(n20345), .ZN(
        n3485) );
  OAI22_X1 U720 ( .A1(n19789), .A2(n18934), .B1(n20620), .B2(n20341), .ZN(
        n3486) );
  OAI22_X1 U721 ( .A1(n19789), .A2(n18935), .B1(n20623), .B2(n20345), .ZN(
        n3487) );
  OAI22_X1 U722 ( .A1(n19789), .A2(n18936), .B1(n20626), .B2(n20344), .ZN(
        n3488) );
  OAI22_X1 U723 ( .A1(n19789), .A2(n18937), .B1(n20629), .B2(n20345), .ZN(
        n3489) );
  OAI22_X1 U724 ( .A1(n19789), .A2(n18938), .B1(n20632), .B2(n20346), .ZN(
        n3490) );
  OAI22_X1 U725 ( .A1(n19790), .A2(n18939), .B1(n20635), .B2(n20346), .ZN(
        n3491) );
  OAI22_X1 U726 ( .A1(n19790), .A2(n18940), .B1(n20638), .B2(n20346), .ZN(
        n3492) );
  OAI22_X1 U727 ( .A1(n19790), .A2(n18941), .B1(n20641), .B2(n20346), .ZN(
        n3493) );
  OAI22_X1 U728 ( .A1(n19790), .A2(n18942), .B1(n20644), .B2(n20346), .ZN(
        n3494) );
  OAI22_X1 U729 ( .A1(n19790), .A2(n18943), .B1(n20647), .B2(n20340), .ZN(
        n3495) );
  OAI22_X1 U730 ( .A1(n19790), .A2(n18944), .B1(n20650), .B2(n20340), .ZN(
        n3496) );
  OAI22_X1 U731 ( .A1(n19790), .A2(n18945), .B1(n20653), .B2(n20340), .ZN(
        n3497) );
  OAI22_X1 U732 ( .A1(n19790), .A2(n18946), .B1(n20656), .B2(n20342), .ZN(
        n3498) );
  OAI22_X1 U733 ( .A1(n19791), .A2(n19395), .B1(n20563), .B2(n20351), .ZN(
        n3499) );
  OAI22_X1 U734 ( .A1(n19791), .A2(n19396), .B1(n20566), .B2(n20349), .ZN(
        n3500) );
  OAI22_X1 U735 ( .A1(n19791), .A2(n19417), .B1(n20569), .B2(n20351), .ZN(
        n3501) );
  OAI22_X1 U736 ( .A1(n19791), .A2(n19397), .B1(n20572), .B2(n20350), .ZN(
        n3502) );
  OAI22_X1 U737 ( .A1(n19791), .A2(n19398), .B1(n20575), .B2(n20349), .ZN(
        n3503) );
  OAI22_X1 U738 ( .A1(n19791), .A2(n19418), .B1(n20578), .B2(n20354), .ZN(
        n3504) );
  OAI22_X1 U739 ( .A1(n19791), .A2(n19399), .B1(n20581), .B2(n20350), .ZN(
        n3505) );
  OAI22_X1 U740 ( .A1(n19791), .A2(n19400), .B1(n20584), .B2(n20351), .ZN(
        n3506) );
  OAI22_X1 U741 ( .A1(n19791), .A2(n19419), .B1(n20587), .B2(n20351), .ZN(
        n3507) );
  OAI22_X1 U742 ( .A1(n19791), .A2(n19401), .B1(n20590), .B2(n20354), .ZN(
        n3508) );
  OAI22_X1 U743 ( .A1(n19791), .A2(n19402), .B1(n20593), .B2(n20352), .ZN(
        n3509) );
  OAI22_X1 U744 ( .A1(n19791), .A2(n19420), .B1(n20596), .B2(n20353), .ZN(
        n3510) );
  OAI22_X1 U745 ( .A1(n19792), .A2(n19403), .B1(n20599), .B2(n20350), .ZN(
        n3511) );
  OAI22_X1 U746 ( .A1(n19792), .A2(n19404), .B1(n20602), .B2(n20351), .ZN(
        n3512) );
  OAI22_X1 U747 ( .A1(n19792), .A2(n19421), .B1(n20605), .B2(n20350), .ZN(
        n3513) );
  OAI22_X1 U748 ( .A1(n19792), .A2(n19405), .B1(n20608), .B2(n20355), .ZN(
        n3514) );
  OAI22_X1 U749 ( .A1(n19792), .A2(n19406), .B1(n20611), .B2(n20352), .ZN(
        n3515) );
  OAI22_X1 U750 ( .A1(n19792), .A2(n19422), .B1(n20614), .B2(n20353), .ZN(
        n3516) );
  OAI22_X1 U751 ( .A1(n19792), .A2(n19407), .B1(n20617), .B2(n20353), .ZN(
        n3517) );
  OAI22_X1 U752 ( .A1(n19792), .A2(n19408), .B1(n20620), .B2(n20349), .ZN(
        n3518) );
  OAI22_X1 U753 ( .A1(n19792), .A2(n19423), .B1(n20623), .B2(n20352), .ZN(
        n3519) );
  OAI22_X1 U754 ( .A1(n19792), .A2(n19409), .B1(n20626), .B2(n20355), .ZN(
        n3520) );
  OAI22_X1 U755 ( .A1(n19792), .A2(n19410), .B1(n20629), .B2(n20355), .ZN(
        n3521) );
  OAI22_X1 U756 ( .A1(n19792), .A2(n19424), .B1(n20632), .B2(n20354), .ZN(
        n3522) );
  OAI22_X1 U757 ( .A1(n19793), .A2(n19411), .B1(n20635), .B2(n20354), .ZN(
        n3523) );
  OAI22_X1 U758 ( .A1(n19793), .A2(n19412), .B1(n20638), .B2(n20355), .ZN(
        n3524) );
  OAI22_X1 U759 ( .A1(n19793), .A2(n19425), .B1(n20641), .B2(n20355), .ZN(
        n3525) );
  OAI22_X1 U760 ( .A1(n19793), .A2(n19413), .B1(n20644), .B2(n20354), .ZN(
        n3526) );
  OAI22_X1 U761 ( .A1(n19793), .A2(n19414), .B1(n20647), .B2(n20351), .ZN(
        n3527) );
  OAI22_X1 U762 ( .A1(n19793), .A2(n19426), .B1(n20650), .B2(n20350), .ZN(
        n3528) );
  OAI22_X1 U763 ( .A1(n19793), .A2(n19415), .B1(n20653), .B2(n20353), .ZN(
        n3529) );
  OAI22_X1 U764 ( .A1(n19793), .A2(n19416), .B1(n20656), .B2(n20352), .ZN(
        n3530) );
  OAI22_X1 U765 ( .A1(n19794), .A2(n18851), .B1(n20563), .B2(n20359), .ZN(
        n3531) );
  OAI22_X1 U766 ( .A1(n19794), .A2(n18852), .B1(n20566), .B2(n20358), .ZN(
        n3532) );
  OAI22_X1 U767 ( .A1(n19794), .A2(n18853), .B1(n20569), .B2(n20359), .ZN(
        n3533) );
  OAI22_X1 U768 ( .A1(n19794), .A2(n18854), .B1(n20572), .B2(n20361), .ZN(
        n3534) );
  OAI22_X1 U769 ( .A1(n19794), .A2(n18855), .B1(n20575), .B2(n20359), .ZN(
        n3535) );
  OAI22_X1 U770 ( .A1(n19794), .A2(n18856), .B1(n20578), .B2(n20364), .ZN(
        n3536) );
  OAI22_X1 U771 ( .A1(n19794), .A2(n18857), .B1(n20581), .B2(n20360), .ZN(
        n3537) );
  OAI22_X1 U772 ( .A1(n19794), .A2(n18858), .B1(n20584), .B2(n20361), .ZN(
        n3538) );
  OAI22_X1 U773 ( .A1(n19794), .A2(n18859), .B1(n20587), .B2(n20361), .ZN(
        n3539) );
  OAI22_X1 U774 ( .A1(n19794), .A2(n18860), .B1(n20590), .B2(n20363), .ZN(
        n3540) );
  OAI22_X1 U775 ( .A1(n19794), .A2(n18861), .B1(n20593), .B2(n20363), .ZN(
        n3541) );
  OAI22_X1 U776 ( .A1(n19794), .A2(n18862), .B1(n20596), .B2(n20362), .ZN(
        n3542) );
  OAI22_X1 U777 ( .A1(n19795), .A2(n18863), .B1(n20599), .B2(n20360), .ZN(
        n3543) );
  OAI22_X1 U778 ( .A1(n19795), .A2(n18864), .B1(n20602), .B2(n20361), .ZN(
        n3544) );
  OAI22_X1 U779 ( .A1(n19795), .A2(n18865), .B1(n20605), .B2(n20360), .ZN(
        n3545) );
  OAI22_X1 U780 ( .A1(n19795), .A2(n18866), .B1(n20608), .B2(n20362), .ZN(
        n3546) );
  OAI22_X1 U781 ( .A1(n19795), .A2(n18867), .B1(n20611), .B2(n20362), .ZN(
        n3547) );
  OAI22_X1 U782 ( .A1(n19795), .A2(n18868), .B1(n20614), .B2(n20362), .ZN(
        n3548) );
  OAI22_X1 U783 ( .A1(n19795), .A2(n18869), .B1(n20617), .B2(n20363), .ZN(
        n3549) );
  OAI22_X1 U784 ( .A1(n19795), .A2(n18870), .B1(n20620), .B2(n20359), .ZN(
        n3550) );
  OAI22_X1 U785 ( .A1(n19795), .A2(n18875), .B1(n20623), .B2(n20363), .ZN(
        n3551) );
  OAI22_X1 U786 ( .A1(n19795), .A2(n18876), .B1(n20626), .B2(n20362), .ZN(
        n3552) );
  OAI22_X1 U787 ( .A1(n19795), .A2(n18877), .B1(n20629), .B2(n20363), .ZN(
        n3553) );
  OAI22_X1 U788 ( .A1(n19795), .A2(n18881), .B1(n20632), .B2(n20364), .ZN(
        n3554) );
  OAI22_X1 U789 ( .A1(n19796), .A2(n18878), .B1(n20635), .B2(n20364), .ZN(
        n3555) );
  OAI22_X1 U790 ( .A1(n19796), .A2(n18879), .B1(n20638), .B2(n20364), .ZN(
        n3556) );
  OAI22_X1 U791 ( .A1(n19796), .A2(n18880), .B1(n20641), .B2(n20364), .ZN(
        n3557) );
  OAI22_X1 U792 ( .A1(n19796), .A2(n18882), .B1(n20644), .B2(n20364), .ZN(
        n3558) );
  OAI22_X1 U793 ( .A1(n19796), .A2(n18871), .B1(n20647), .B2(n20358), .ZN(
        n3559) );
  OAI22_X1 U794 ( .A1(n19796), .A2(n18872), .B1(n20650), .B2(n20358), .ZN(
        n3560) );
  OAI22_X1 U795 ( .A1(n19796), .A2(n18873), .B1(n20653), .B2(n20358), .ZN(
        n3561) );
  OAI22_X1 U796 ( .A1(n19796), .A2(n18874), .B1(n20656), .B2(n20360), .ZN(
        n3562) );
  OAI22_X1 U797 ( .A1(n19782), .A2(n19332), .B1(n20561), .B2(n20324), .ZN(
        n3279) );
  OAI22_X1 U798 ( .A1(n19782), .A2(n19355), .B1(n20564), .B2(n20322), .ZN(
        n3284) );
  OAI22_X1 U799 ( .A1(n19782), .A2(n19333), .B1(n20567), .B2(n20324), .ZN(
        n3289) );
  OAI22_X1 U800 ( .A1(n19782), .A2(n19334), .B1(n20570), .B2(n20323), .ZN(
        n3294) );
  OAI22_X1 U801 ( .A1(n19782), .A2(n19335), .B1(n20573), .B2(n20322), .ZN(
        n3299) );
  OAI22_X1 U802 ( .A1(n19782), .A2(n19356), .B1(n20576), .B2(n20327), .ZN(
        n3304) );
  OAI22_X1 U803 ( .A1(n19782), .A2(n19336), .B1(n20579), .B2(n20323), .ZN(
        n3309) );
  OAI22_X1 U804 ( .A1(n19782), .A2(n19337), .B1(n20582), .B2(n20324), .ZN(
        n3314) );
  OAI22_X1 U805 ( .A1(n19782), .A2(n19338), .B1(n20585), .B2(n20324), .ZN(
        n3319) );
  OAI22_X1 U806 ( .A1(n19782), .A2(n19357), .B1(n20588), .B2(n20327), .ZN(
        n3324) );
  OAI22_X1 U807 ( .A1(n19782), .A2(n19339), .B1(n20591), .B2(n20325), .ZN(
        n3329) );
  OAI22_X1 U808 ( .A1(n19782), .A2(n19340), .B1(n20594), .B2(n20326), .ZN(
        n3334) );
  OAI22_X1 U809 ( .A1(n19783), .A2(n19358), .B1(n20597), .B2(n20323), .ZN(
        n3339) );
  OAI22_X1 U810 ( .A1(n19783), .A2(n19341), .B1(n20600), .B2(n20324), .ZN(
        n3344) );
  OAI22_X1 U811 ( .A1(n19783), .A2(n19342), .B1(n20603), .B2(n20323), .ZN(
        n3349) );
  OAI22_X1 U812 ( .A1(n19783), .A2(n19343), .B1(n20606), .B2(n20328), .ZN(
        n3354) );
  OAI22_X1 U813 ( .A1(n19783), .A2(n19359), .B1(n20609), .B2(n20325), .ZN(
        n3359) );
  OAI22_X1 U814 ( .A1(n19783), .A2(n19344), .B1(n20612), .B2(n20326), .ZN(
        n3364) );
  OAI22_X1 U815 ( .A1(n19783), .A2(n19345), .B1(n20615), .B2(n20326), .ZN(
        n3369) );
  OAI22_X1 U816 ( .A1(n19783), .A2(n19346), .B1(n20618), .B2(n20322), .ZN(
        n3374) );
  OAI22_X1 U817 ( .A1(n19783), .A2(n19347), .B1(n20621), .B2(n20325), .ZN(
        n3379) );
  OAI22_X1 U818 ( .A1(n19783), .A2(n19348), .B1(n20624), .B2(n20328), .ZN(
        n3384) );
  OAI22_X1 U819 ( .A1(n19783), .A2(n19349), .B1(n20627), .B2(n20328), .ZN(
        n3389) );
  OAI22_X1 U820 ( .A1(n19783), .A2(n19360), .B1(n20630), .B2(n20327), .ZN(
        n3394) );
  OAI22_X1 U821 ( .A1(n19784), .A2(n19350), .B1(n20633), .B2(n20327), .ZN(
        n3399) );
  OAI22_X1 U822 ( .A1(n19784), .A2(n19351), .B1(n20636), .B2(n20328), .ZN(
        n3404) );
  OAI22_X1 U823 ( .A1(n19784), .A2(n19352), .B1(n20639), .B2(n20328), .ZN(
        n3409) );
  OAI22_X1 U824 ( .A1(n19784), .A2(n19361), .B1(n20642), .B2(n20327), .ZN(
        n3414) );
  OAI22_X1 U825 ( .A1(n19784), .A2(n19353), .B1(n20645), .B2(n20324), .ZN(
        n3419) );
  OAI22_X1 U826 ( .A1(n19784), .A2(n19354), .B1(n20648), .B2(n20323), .ZN(
        n3424) );
  OAI22_X1 U827 ( .A1(n19784), .A2(n19362), .B1(n20651), .B2(n20326), .ZN(
        n3429) );
  OAI22_X1 U828 ( .A1(n19784), .A2(n19331), .B1(n20654), .B2(n20325), .ZN(
        n3434) );
  OAI22_X1 U829 ( .A1(n19806), .A2(n19267), .B1(n20562), .B2(n20396), .ZN(
        n3659) );
  OAI22_X1 U830 ( .A1(n19806), .A2(n19268), .B1(n20565), .B2(n20394), .ZN(
        n3660) );
  OAI22_X1 U831 ( .A1(n19806), .A2(n19269), .B1(n20568), .B2(n20396), .ZN(
        n3661) );
  OAI22_X1 U832 ( .A1(n19806), .A2(n19270), .B1(n20571), .B2(n20395), .ZN(
        n3662) );
  OAI22_X1 U833 ( .A1(n19806), .A2(n19271), .B1(n20574), .B2(n20394), .ZN(
        n3663) );
  OAI22_X1 U834 ( .A1(n19806), .A2(n19272), .B1(n20577), .B2(n20399), .ZN(
        n3664) );
  OAI22_X1 U835 ( .A1(n19806), .A2(n19273), .B1(n20580), .B2(n20395), .ZN(
        n3665) );
  OAI22_X1 U836 ( .A1(n19806), .A2(n19274), .B1(n20583), .B2(n20396), .ZN(
        n3666) );
  OAI22_X1 U837 ( .A1(n19806), .A2(n19275), .B1(n20586), .B2(n20396), .ZN(
        n3667) );
  OAI22_X1 U838 ( .A1(n19806), .A2(n19276), .B1(n20589), .B2(n20399), .ZN(
        n3668) );
  OAI22_X1 U839 ( .A1(n19806), .A2(n19277), .B1(n20592), .B2(n20397), .ZN(
        n3669) );
  OAI22_X1 U840 ( .A1(n19806), .A2(n19278), .B1(n20595), .B2(n20398), .ZN(
        n3670) );
  OAI22_X1 U841 ( .A1(n19807), .A2(n19279), .B1(n20598), .B2(n20395), .ZN(
        n3671) );
  OAI22_X1 U842 ( .A1(n19807), .A2(n19280), .B1(n20601), .B2(n20396), .ZN(
        n3672) );
  OAI22_X1 U843 ( .A1(n19807), .A2(n19281), .B1(n20604), .B2(n20395), .ZN(
        n3673) );
  OAI22_X1 U844 ( .A1(n19807), .A2(n19282), .B1(n20607), .B2(n20400), .ZN(
        n3674) );
  OAI22_X1 U845 ( .A1(n19807), .A2(n19283), .B1(n20610), .B2(n20397), .ZN(
        n3675) );
  OAI22_X1 U846 ( .A1(n19807), .A2(n19284), .B1(n20613), .B2(n20398), .ZN(
        n3676) );
  OAI22_X1 U847 ( .A1(n19807), .A2(n19285), .B1(n20616), .B2(n20398), .ZN(
        n3677) );
  OAI22_X1 U848 ( .A1(n19807), .A2(n19286), .B1(n20619), .B2(n20394), .ZN(
        n3678) );
  OAI22_X1 U849 ( .A1(n19807), .A2(n19287), .B1(n20622), .B2(n20397), .ZN(
        n3679) );
  OAI22_X1 U850 ( .A1(n19807), .A2(n19288), .B1(n20625), .B2(n20400), .ZN(
        n3680) );
  OAI22_X1 U851 ( .A1(n19807), .A2(n19289), .B1(n20628), .B2(n20400), .ZN(
        n3681) );
  OAI22_X1 U852 ( .A1(n19807), .A2(n19290), .B1(n20631), .B2(n20399), .ZN(
        n3682) );
  OAI22_X1 U853 ( .A1(n19808), .A2(n19291), .B1(n20634), .B2(n20399), .ZN(
        n3683) );
  OAI22_X1 U854 ( .A1(n19808), .A2(n19292), .B1(n20637), .B2(n20400), .ZN(
        n3684) );
  OAI22_X1 U855 ( .A1(n19808), .A2(n19293), .B1(n20640), .B2(n20400), .ZN(
        n3685) );
  OAI22_X1 U856 ( .A1(n19808), .A2(n19294), .B1(n20643), .B2(n20399), .ZN(
        n3686) );
  OAI22_X1 U857 ( .A1(n19808), .A2(n19295), .B1(n20646), .B2(n20396), .ZN(
        n3687) );
  OAI22_X1 U858 ( .A1(n19808), .A2(n19296), .B1(n20649), .B2(n20395), .ZN(
        n3688) );
  OAI22_X1 U859 ( .A1(n19808), .A2(n19297), .B1(n20652), .B2(n20398), .ZN(
        n3689) );
  OAI22_X1 U860 ( .A1(n19808), .A2(n19298), .B1(n20655), .B2(n20397), .ZN(
        n3690) );
  OAI22_X1 U861 ( .A1(n19809), .A2(n18883), .B1(n20562), .B2(n20404), .ZN(
        n3691) );
  OAI22_X1 U862 ( .A1(n19809), .A2(n18884), .B1(n20565), .B2(n20403), .ZN(
        n3692) );
  OAI22_X1 U863 ( .A1(n19809), .A2(n18885), .B1(n20568), .B2(n20404), .ZN(
        n3693) );
  OAI22_X1 U864 ( .A1(n19809), .A2(n18886), .B1(n20571), .B2(n20406), .ZN(
        n3694) );
  OAI22_X1 U865 ( .A1(n19809), .A2(n18887), .B1(n20574), .B2(n20404), .ZN(
        n3695) );
  OAI22_X1 U866 ( .A1(n19809), .A2(n18888), .B1(n20577), .B2(n20409), .ZN(
        n3696) );
  OAI22_X1 U867 ( .A1(n19809), .A2(n18889), .B1(n20580), .B2(n20405), .ZN(
        n3697) );
  OAI22_X1 U868 ( .A1(n19809), .A2(n18890), .B1(n20583), .B2(n20406), .ZN(
        n3698) );
  OAI22_X1 U869 ( .A1(n19809), .A2(n18891), .B1(n20586), .B2(n20406), .ZN(
        n3699) );
  OAI22_X1 U870 ( .A1(n19809), .A2(n18892), .B1(n20589), .B2(n20408), .ZN(
        n3700) );
  OAI22_X1 U871 ( .A1(n19809), .A2(n18893), .B1(n20592), .B2(n20408), .ZN(
        n3701) );
  OAI22_X1 U872 ( .A1(n19809), .A2(n18894), .B1(n20595), .B2(n20407), .ZN(
        n3702) );
  OAI22_X1 U873 ( .A1(n19810), .A2(n18895), .B1(n20598), .B2(n20405), .ZN(
        n3703) );
  OAI22_X1 U874 ( .A1(n19810), .A2(n18896), .B1(n20601), .B2(n20406), .ZN(
        n3704) );
  OAI22_X1 U875 ( .A1(n19810), .A2(n18897), .B1(n20604), .B2(n20405), .ZN(
        n3705) );
  OAI22_X1 U876 ( .A1(n19810), .A2(n18898), .B1(n20607), .B2(n20407), .ZN(
        n3706) );
  OAI22_X1 U877 ( .A1(n19810), .A2(n18899), .B1(n20610), .B2(n20407), .ZN(
        n3707) );
  OAI22_X1 U878 ( .A1(n19810), .A2(n18900), .B1(n20613), .B2(n20407), .ZN(
        n3708) );
  OAI22_X1 U879 ( .A1(n19810), .A2(n18901), .B1(n20616), .B2(n20408), .ZN(
        n3709) );
  OAI22_X1 U880 ( .A1(n19810), .A2(n18902), .B1(n20619), .B2(n20404), .ZN(
        n3710) );
  OAI22_X1 U881 ( .A1(n19810), .A2(n18907), .B1(n20622), .B2(n20408), .ZN(
        n3711) );
  OAI22_X1 U882 ( .A1(n19810), .A2(n18908), .B1(n20625), .B2(n20407), .ZN(
        n3712) );
  OAI22_X1 U883 ( .A1(n19810), .A2(n18909), .B1(n20628), .B2(n20408), .ZN(
        n3713) );
  OAI22_X1 U884 ( .A1(n19810), .A2(n18910), .B1(n20631), .B2(n20409), .ZN(
        n3714) );
  OAI22_X1 U885 ( .A1(n19811), .A2(n18911), .B1(n20634), .B2(n20409), .ZN(
        n3715) );
  OAI22_X1 U886 ( .A1(n19811), .A2(n18912), .B1(n20637), .B2(n20409), .ZN(
        n3716) );
  OAI22_X1 U887 ( .A1(n19811), .A2(n18913), .B1(n20640), .B2(n20409), .ZN(
        n3717) );
  OAI22_X1 U888 ( .A1(n19811), .A2(n18914), .B1(n20643), .B2(n20409), .ZN(
        n3718) );
  OAI22_X1 U889 ( .A1(n19811), .A2(n18903), .B1(n20646), .B2(n20403), .ZN(
        n3719) );
  OAI22_X1 U890 ( .A1(n19811), .A2(n18904), .B1(n20649), .B2(n20403), .ZN(
        n3720) );
  OAI22_X1 U891 ( .A1(n19811), .A2(n18905), .B1(n20652), .B2(n20403), .ZN(
        n3721) );
  OAI22_X1 U892 ( .A1(n19811), .A2(n18906), .B1(n20655), .B2(n20405), .ZN(
        n3722) );
  OAI22_X1 U893 ( .A1(n19812), .A2(n19043), .B1(n20562), .B2(n20414), .ZN(
        n3723) );
  OAI22_X1 U894 ( .A1(n19812), .A2(n19044), .B1(n20565), .B2(n20412), .ZN(
        n3724) );
  OAI22_X1 U895 ( .A1(n19812), .A2(n19045), .B1(n20568), .B2(n20414), .ZN(
        n3725) );
  OAI22_X1 U896 ( .A1(n19812), .A2(n19046), .B1(n20571), .B2(n20413), .ZN(
        n3726) );
  OAI22_X1 U897 ( .A1(n19812), .A2(n19047), .B1(n20574), .B2(n20412), .ZN(
        n3727) );
  OAI22_X1 U898 ( .A1(n19812), .A2(n19048), .B1(n20577), .B2(n20417), .ZN(
        n3728) );
  OAI22_X1 U899 ( .A1(n19812), .A2(n19049), .B1(n20580), .B2(n20413), .ZN(
        n3729) );
  OAI22_X1 U900 ( .A1(n19812), .A2(n19050), .B1(n20583), .B2(n20414), .ZN(
        n3730) );
  OAI22_X1 U901 ( .A1(n19812), .A2(n19051), .B1(n20586), .B2(n20414), .ZN(
        n3731) );
  OAI22_X1 U902 ( .A1(n19812), .A2(n19052), .B1(n20589), .B2(n20417), .ZN(
        n3732) );
  OAI22_X1 U903 ( .A1(n19812), .A2(n19053), .B1(n20592), .B2(n20415), .ZN(
        n3733) );
  OAI22_X1 U904 ( .A1(n19812), .A2(n19054), .B1(n20595), .B2(n20416), .ZN(
        n3734) );
  OAI22_X1 U905 ( .A1(n19813), .A2(n19055), .B1(n20598), .B2(n20413), .ZN(
        n3735) );
  OAI22_X1 U906 ( .A1(n19813), .A2(n19056), .B1(n20601), .B2(n20414), .ZN(
        n3736) );
  OAI22_X1 U907 ( .A1(n19813), .A2(n19057), .B1(n20604), .B2(n20413), .ZN(
        n3737) );
  OAI22_X1 U908 ( .A1(n19813), .A2(n19058), .B1(n20607), .B2(n20418), .ZN(
        n3738) );
  OAI22_X1 U909 ( .A1(n19813), .A2(n19059), .B1(n20610), .B2(n20415), .ZN(
        n3739) );
  OAI22_X1 U910 ( .A1(n19813), .A2(n19060), .B1(n20613), .B2(n20416), .ZN(
        n3740) );
  OAI22_X1 U911 ( .A1(n19813), .A2(n19061), .B1(n20616), .B2(n20416), .ZN(
        n3741) );
  OAI22_X1 U912 ( .A1(n19813), .A2(n19062), .B1(n20619), .B2(n20412), .ZN(
        n3742) );
  OAI22_X1 U913 ( .A1(n19813), .A2(n19063), .B1(n20622), .B2(n20415), .ZN(
        n3743) );
  OAI22_X1 U914 ( .A1(n19813), .A2(n19064), .B1(n20625), .B2(n20418), .ZN(
        n3744) );
  OAI22_X1 U915 ( .A1(n19813), .A2(n19065), .B1(n20628), .B2(n20418), .ZN(
        n3745) );
  OAI22_X1 U916 ( .A1(n19813), .A2(n19066), .B1(n20631), .B2(n20417), .ZN(
        n3746) );
  OAI22_X1 U917 ( .A1(n19814), .A2(n19067), .B1(n20634), .B2(n20417), .ZN(
        n3747) );
  OAI22_X1 U918 ( .A1(n19814), .A2(n19068), .B1(n20637), .B2(n20418), .ZN(
        n3748) );
  OAI22_X1 U919 ( .A1(n19814), .A2(n19069), .B1(n20640), .B2(n20418), .ZN(
        n3749) );
  OAI22_X1 U920 ( .A1(n19814), .A2(n19070), .B1(n20643), .B2(n20417), .ZN(
        n3750) );
  OAI22_X1 U921 ( .A1(n19814), .A2(n19071), .B1(n20646), .B2(n20414), .ZN(
        n3751) );
  OAI22_X1 U922 ( .A1(n19814), .A2(n19072), .B1(n20649), .B2(n20413), .ZN(
        n3752) );
  OAI22_X1 U923 ( .A1(n19814), .A2(n19073), .B1(n20652), .B2(n20416), .ZN(
        n3753) );
  OAI22_X1 U924 ( .A1(n19814), .A2(n19074), .B1(n20655), .B2(n20415), .ZN(
        n3754) );
  OAI22_X1 U925 ( .A1(n19818), .A2(n19235), .B1(n20562), .B2(n20432), .ZN(
        n3787) );
  OAI22_X1 U926 ( .A1(n19818), .A2(n19236), .B1(n20565), .B2(n20430), .ZN(
        n3788) );
  OAI22_X1 U927 ( .A1(n19818), .A2(n19237), .B1(n20568), .B2(n20432), .ZN(
        n3789) );
  OAI22_X1 U928 ( .A1(n19818), .A2(n19238), .B1(n20571), .B2(n20431), .ZN(
        n3790) );
  OAI22_X1 U929 ( .A1(n19818), .A2(n19239), .B1(n20574), .B2(n20430), .ZN(
        n3791) );
  OAI22_X1 U930 ( .A1(n19818), .A2(n19240), .B1(n20577), .B2(n20435), .ZN(
        n3792) );
  OAI22_X1 U931 ( .A1(n19818), .A2(n19241), .B1(n20580), .B2(n20431), .ZN(
        n3793) );
  OAI22_X1 U932 ( .A1(n19818), .A2(n19242), .B1(n20583), .B2(n20432), .ZN(
        n3794) );
  OAI22_X1 U933 ( .A1(n19818), .A2(n19243), .B1(n20586), .B2(n20432), .ZN(
        n3795) );
  OAI22_X1 U934 ( .A1(n19818), .A2(n19244), .B1(n20589), .B2(n20435), .ZN(
        n3796) );
  OAI22_X1 U935 ( .A1(n19818), .A2(n19245), .B1(n20592), .B2(n20433), .ZN(
        n3797) );
  OAI22_X1 U936 ( .A1(n19818), .A2(n19246), .B1(n20595), .B2(n20434), .ZN(
        n3798) );
  OAI22_X1 U937 ( .A1(n19819), .A2(n19247), .B1(n20598), .B2(n20431), .ZN(
        n3799) );
  OAI22_X1 U938 ( .A1(n19819), .A2(n19248), .B1(n20601), .B2(n20432), .ZN(
        n3800) );
  OAI22_X1 U939 ( .A1(n19819), .A2(n19249), .B1(n20604), .B2(n20431), .ZN(
        n3801) );
  OAI22_X1 U940 ( .A1(n19819), .A2(n19250), .B1(n20607), .B2(n20436), .ZN(
        n3802) );
  OAI22_X1 U941 ( .A1(n19819), .A2(n19251), .B1(n20610), .B2(n20433), .ZN(
        n3803) );
  OAI22_X1 U942 ( .A1(n19819), .A2(n19252), .B1(n20613), .B2(n20434), .ZN(
        n3804) );
  OAI22_X1 U943 ( .A1(n19819), .A2(n19253), .B1(n20616), .B2(n20434), .ZN(
        n3805) );
  OAI22_X1 U944 ( .A1(n19819), .A2(n19254), .B1(n20619), .B2(n20430), .ZN(
        n3806) );
  OAI22_X1 U945 ( .A1(n19819), .A2(n19259), .B1(n20622), .B2(n20433), .ZN(
        n3807) );
  OAI22_X1 U946 ( .A1(n19819), .A2(n19260), .B1(n20625), .B2(n20436), .ZN(
        n3808) );
  OAI22_X1 U947 ( .A1(n19819), .A2(n19261), .B1(n20628), .B2(n20436), .ZN(
        n3809) );
  OAI22_X1 U948 ( .A1(n19819), .A2(n19265), .B1(n20631), .B2(n20435), .ZN(
        n3810) );
  OAI22_X1 U949 ( .A1(n19820), .A2(n19262), .B1(n20634), .B2(n20435), .ZN(
        n3811) );
  OAI22_X1 U950 ( .A1(n19820), .A2(n19263), .B1(n20637), .B2(n20436), .ZN(
        n3812) );
  OAI22_X1 U951 ( .A1(n19820), .A2(n19264), .B1(n20640), .B2(n20436), .ZN(
        n3813) );
  OAI22_X1 U952 ( .A1(n19820), .A2(n19266), .B1(n20643), .B2(n20435), .ZN(
        n3814) );
  OAI22_X1 U953 ( .A1(n19820), .A2(n19255), .B1(n20646), .B2(n20432), .ZN(
        n3815) );
  OAI22_X1 U954 ( .A1(n19820), .A2(n19256), .B1(n20649), .B2(n20431), .ZN(
        n3816) );
  OAI22_X1 U955 ( .A1(n19820), .A2(n19257), .B1(n20652), .B2(n20434), .ZN(
        n3817) );
  OAI22_X1 U956 ( .A1(n19820), .A2(n19258), .B1(n20655), .B2(n20433), .ZN(
        n3818) );
  OAI22_X1 U957 ( .A1(n19821), .A2(n19107), .B1(n20562), .B2(n20441), .ZN(
        n3819) );
  OAI22_X1 U958 ( .A1(n19821), .A2(n19108), .B1(n20565), .B2(n20439), .ZN(
        n3820) );
  OAI22_X1 U959 ( .A1(n19821), .A2(n19109), .B1(n20568), .B2(n20441), .ZN(
        n3821) );
  OAI22_X1 U960 ( .A1(n19821), .A2(n19110), .B1(n20571), .B2(n20440), .ZN(
        n3822) );
  OAI22_X1 U961 ( .A1(n19821), .A2(n19111), .B1(n20574), .B2(n20439), .ZN(
        n3823) );
  OAI22_X1 U962 ( .A1(n19821), .A2(n19112), .B1(n20577), .B2(n20444), .ZN(
        n3824) );
  OAI22_X1 U963 ( .A1(n19821), .A2(n19113), .B1(n20580), .B2(n20440), .ZN(
        n3825) );
  OAI22_X1 U964 ( .A1(n19821), .A2(n19114), .B1(n20583), .B2(n20441), .ZN(
        n3826) );
  OAI22_X1 U965 ( .A1(n19821), .A2(n19115), .B1(n20586), .B2(n20441), .ZN(
        n3827) );
  OAI22_X1 U966 ( .A1(n19821), .A2(n19116), .B1(n20589), .B2(n20444), .ZN(
        n3828) );
  OAI22_X1 U967 ( .A1(n19821), .A2(n19117), .B1(n20592), .B2(n20442), .ZN(
        n3829) );
  OAI22_X1 U968 ( .A1(n19821), .A2(n19118), .B1(n20595), .B2(n20443), .ZN(
        n3830) );
  OAI22_X1 U969 ( .A1(n19822), .A2(n19119), .B1(n20598), .B2(n20440), .ZN(
        n3831) );
  OAI22_X1 U970 ( .A1(n19822), .A2(n19120), .B1(n20601), .B2(n20441), .ZN(
        n3832) );
  OAI22_X1 U971 ( .A1(n19822), .A2(n19121), .B1(n20604), .B2(n20440), .ZN(
        n3833) );
  OAI22_X1 U972 ( .A1(n19822), .A2(n19122), .B1(n20607), .B2(n20445), .ZN(
        n3834) );
  OAI22_X1 U973 ( .A1(n19822), .A2(n19123), .B1(n20610), .B2(n20442), .ZN(
        n3835) );
  OAI22_X1 U974 ( .A1(n19822), .A2(n19124), .B1(n20613), .B2(n20443), .ZN(
        n3836) );
  OAI22_X1 U975 ( .A1(n19822), .A2(n19125), .B1(n20616), .B2(n20443), .ZN(
        n3837) );
  OAI22_X1 U976 ( .A1(n19822), .A2(n19126), .B1(n20619), .B2(n20439), .ZN(
        n3838) );
  OAI22_X1 U977 ( .A1(n19822), .A2(n19127), .B1(n20622), .B2(n20442), .ZN(
        n3839) );
  OAI22_X1 U978 ( .A1(n19822), .A2(n19128), .B1(n20625), .B2(n20445), .ZN(
        n3840) );
  OAI22_X1 U979 ( .A1(n19822), .A2(n19129), .B1(n20628), .B2(n20445), .ZN(
        n3841) );
  OAI22_X1 U980 ( .A1(n19822), .A2(n19130), .B1(n20631), .B2(n20444), .ZN(
        n3842) );
  OAI22_X1 U981 ( .A1(n19823), .A2(n19131), .B1(n20634), .B2(n20444), .ZN(
        n3843) );
  OAI22_X1 U982 ( .A1(n19823), .A2(n19132), .B1(n20637), .B2(n20445), .ZN(
        n3844) );
  OAI22_X1 U983 ( .A1(n19823), .A2(n19133), .B1(n20640), .B2(n20445), .ZN(
        n3845) );
  OAI22_X1 U984 ( .A1(n19823), .A2(n19134), .B1(n20643), .B2(n20444), .ZN(
        n3846) );
  OAI22_X1 U985 ( .A1(n19823), .A2(n19135), .B1(n20646), .B2(n20441), .ZN(
        n3847) );
  OAI22_X1 U986 ( .A1(n19823), .A2(n19136), .B1(n20649), .B2(n20440), .ZN(
        n3848) );
  OAI22_X1 U987 ( .A1(n19823), .A2(n19137), .B1(n20652), .B2(n20443), .ZN(
        n3849) );
  OAI22_X1 U988 ( .A1(n19823), .A2(n19138), .B1(n20655), .B2(n20442), .ZN(
        n3850) );
  OAI22_X1 U989 ( .A1(n19833), .A2(n19427), .B1(n20561), .B2(n20474), .ZN(
        n3947) );
  OAI22_X1 U990 ( .A1(n19833), .A2(n19443), .B1(n20564), .B2(n20475), .ZN(
        n3948) );
  OAI22_X1 U991 ( .A1(n19833), .A2(n19449), .B1(n20567), .B2(n20474), .ZN(
        n3949) );
  OAI22_X1 U992 ( .A1(n19833), .A2(n19428), .B1(n20570), .B2(n20475), .ZN(
        n3950) );
  OAI22_X1 U993 ( .A1(n19833), .A2(n19429), .B1(n20573), .B2(n20476), .ZN(
        n3951) );
  OAI22_X1 U994 ( .A1(n19833), .A2(n19457), .B1(n20576), .B2(n20474), .ZN(
        n3952) );
  OAI22_X1 U995 ( .A1(n19833), .A2(n19430), .B1(n20579), .B2(n20476), .ZN(
        n3953) );
  OAI22_X1 U996 ( .A1(n19833), .A2(n19431), .B1(n20582), .B2(n20477), .ZN(
        n3954) );
  OAI22_X1 U997 ( .A1(n19833), .A2(n19450), .B1(n20585), .B2(n20477), .ZN(
        n3955) );
  OAI22_X1 U998 ( .A1(n19833), .A2(n19444), .B1(n20588), .B2(n20478), .ZN(
        n3956) );
  OAI22_X1 U999 ( .A1(n19833), .A2(n19432), .B1(n20591), .B2(n20479), .ZN(
        n3957) );
  OAI22_X1 U1000 ( .A1(n19833), .A2(n19451), .B1(n20594), .B2(n20475), .ZN(
        n3958) );
  OAI22_X1 U1001 ( .A1(n19834), .A2(n19445), .B1(n20597), .B2(n20478), .ZN(
        n3959) );
  OAI22_X1 U1002 ( .A1(n19834), .A2(n19433), .B1(n20600), .B2(n20479), .ZN(
        n3960) );
  OAI22_X1 U1003 ( .A1(n19834), .A2(n19452), .B1(n20603), .B2(n20474), .ZN(
        n3961) );
  OAI22_X1 U1004 ( .A1(n19834), .A2(n19434), .B1(n20606), .B2(n20475), .ZN(
        n3962) );
  OAI22_X1 U1005 ( .A1(n19834), .A2(n19446), .B1(n20609), .B2(n20476), .ZN(
        n3963) );
  OAI22_X1 U1006 ( .A1(n19834), .A2(n19453), .B1(n20612), .B2(n20476), .ZN(
        n3964) );
  OAI22_X1 U1007 ( .A1(n19834), .A2(n19435), .B1(n20615), .B2(n20474), .ZN(
        n3965) );
  OAI22_X1 U1008 ( .A1(n19834), .A2(n19436), .B1(n20618), .B2(n20475), .ZN(
        n3966) );
  OAI22_X1 U1009 ( .A1(n19834), .A2(n19454), .B1(n20621), .B2(n20477), .ZN(
        n3967) );
  OAI22_X1 U1010 ( .A1(n19834), .A2(n19437), .B1(n20624), .B2(n20478), .ZN(
        n3968) );
  OAI22_X1 U1011 ( .A1(n19834), .A2(n19438), .B1(n20627), .B2(n20479), .ZN(
        n3969) );
  OAI22_X1 U1012 ( .A1(n19834), .A2(n19458), .B1(n20630), .B2(n20477), .ZN(
        n3970) );
  OAI22_X1 U1013 ( .A1(n19835), .A2(n19439), .B1(n20633), .B2(n20476), .ZN(
        n3971) );
  OAI22_X1 U1014 ( .A1(n19835), .A2(n19440), .B1(n20636), .B2(n20477), .ZN(
        n3972) );
  OAI22_X1 U1015 ( .A1(n19835), .A2(n19455), .B1(n20639), .B2(n20474), .ZN(
        n3973) );
  OAI22_X1 U1016 ( .A1(n19835), .A2(n19447), .B1(n20642), .B2(n20475), .ZN(
        n3974) );
  OAI22_X1 U1017 ( .A1(n19835), .A2(n19441), .B1(n20645), .B2(n20476), .ZN(
        n3975) );
  OAI22_X1 U1018 ( .A1(n19835), .A2(n19456), .B1(n20648), .B2(n20478), .ZN(
        n3976) );
  OAI22_X1 U1019 ( .A1(n19835), .A2(n19448), .B1(n20651), .B2(n20478), .ZN(
        n3977) );
  OAI22_X1 U1020 ( .A1(n19835), .A2(n19442), .B1(n20654), .B2(n20479), .ZN(
        n3978) );
  OAI22_X1 U1021 ( .A1(n19836), .A2(n19299), .B1(n20561), .B2(n20484), .ZN(
        n3979) );
  OAI22_X1 U1022 ( .A1(n19836), .A2(n19300), .B1(n20564), .B2(n20482), .ZN(
        n3980) );
  OAI22_X1 U1023 ( .A1(n19836), .A2(n19321), .B1(n20567), .B2(n20484), .ZN(
        n3981) );
  OAI22_X1 U1024 ( .A1(n19836), .A2(n19301), .B1(n20570), .B2(n20483), .ZN(
        n3982) );
  OAI22_X1 U1025 ( .A1(n19836), .A2(n19302), .B1(n20573), .B2(n20482), .ZN(
        n3983) );
  OAI22_X1 U1026 ( .A1(n19836), .A2(n19322), .B1(n20576), .B2(n20487), .ZN(
        n3984) );
  OAI22_X1 U1027 ( .A1(n19836), .A2(n19303), .B1(n20579), .B2(n20483), .ZN(
        n3985) );
  OAI22_X1 U1028 ( .A1(n19836), .A2(n19304), .B1(n20582), .B2(n20484), .ZN(
        n3986) );
  OAI22_X1 U1029 ( .A1(n19836), .A2(n19323), .B1(n20585), .B2(n20484), .ZN(
        n3987) );
  OAI22_X1 U1030 ( .A1(n19836), .A2(n19305), .B1(n20588), .B2(n20487), .ZN(
        n3988) );
  OAI22_X1 U1031 ( .A1(n19836), .A2(n19306), .B1(n20591), .B2(n20485), .ZN(
        n3989) );
  OAI22_X1 U1032 ( .A1(n19836), .A2(n19324), .B1(n20594), .B2(n20486), .ZN(
        n3990) );
  OAI22_X1 U1033 ( .A1(n19837), .A2(n19307), .B1(n20597), .B2(n20483), .ZN(
        n3991) );
  OAI22_X1 U1034 ( .A1(n19837), .A2(n19308), .B1(n20600), .B2(n20484), .ZN(
        n3992) );
  OAI22_X1 U1035 ( .A1(n19837), .A2(n19325), .B1(n20603), .B2(n20483), .ZN(
        n3993) );
  OAI22_X1 U1036 ( .A1(n19837), .A2(n19309), .B1(n20606), .B2(n20488), .ZN(
        n3994) );
  OAI22_X1 U1037 ( .A1(n19837), .A2(n19310), .B1(n20609), .B2(n20485), .ZN(
        n3995) );
  OAI22_X1 U1038 ( .A1(n19837), .A2(n19326), .B1(n20612), .B2(n20486), .ZN(
        n3996) );
  OAI22_X1 U1039 ( .A1(n19837), .A2(n19311), .B1(n20615), .B2(n20486), .ZN(
        n3997) );
  OAI22_X1 U1040 ( .A1(n19837), .A2(n19312), .B1(n20618), .B2(n20482), .ZN(
        n3998) );
  OAI22_X1 U1041 ( .A1(n19837), .A2(n19327), .B1(n20621), .B2(n20485), .ZN(
        n3999) );
  OAI22_X1 U1042 ( .A1(n19837), .A2(n19313), .B1(n20624), .B2(n20488), .ZN(
        n4000) );
  OAI22_X1 U1043 ( .A1(n19837), .A2(n19314), .B1(n20627), .B2(n20488), .ZN(
        n4001) );
  OAI22_X1 U1044 ( .A1(n19837), .A2(n19328), .B1(n20630), .B2(n20487), .ZN(
        n4002) );
  OAI22_X1 U1045 ( .A1(n19838), .A2(n19315), .B1(n20633), .B2(n20487), .ZN(
        n4003) );
  OAI22_X1 U1046 ( .A1(n19838), .A2(n19316), .B1(n20636), .B2(n20488), .ZN(
        n4004) );
  OAI22_X1 U1047 ( .A1(n19838), .A2(n19329), .B1(n20639), .B2(n20488), .ZN(
        n4005) );
  OAI22_X1 U1048 ( .A1(n19838), .A2(n19317), .B1(n20642), .B2(n20487), .ZN(
        n4006) );
  OAI22_X1 U1049 ( .A1(n19838), .A2(n19318), .B1(n20645), .B2(n20484), .ZN(
        n4007) );
  OAI22_X1 U1050 ( .A1(n19838), .A2(n19330), .B1(n20648), .B2(n20483), .ZN(
        n4008) );
  OAI22_X1 U1051 ( .A1(n19838), .A2(n19319), .B1(n20651), .B2(n20486), .ZN(
        n4009) );
  OAI22_X1 U1052 ( .A1(n19838), .A2(n19320), .B1(n20654), .B2(n20485), .ZN(
        n4010) );
  OAI22_X1 U1053 ( .A1(n19845), .A2(n18947), .B1(n20561), .B2(n20508), .ZN(
        n4075) );
  OAI22_X1 U1054 ( .A1(n19845), .A2(n18948), .B1(n20564), .B2(n20507), .ZN(
        n4076) );
  OAI22_X1 U1055 ( .A1(n19845), .A2(n18949), .B1(n20567), .B2(n20508), .ZN(
        n4077) );
  OAI22_X1 U1056 ( .A1(n19845), .A2(n18950), .B1(n20570), .B2(n20510), .ZN(
        n4078) );
  OAI22_X1 U1057 ( .A1(n19845), .A2(n18951), .B1(n20573), .B2(n20508), .ZN(
        n4079) );
  OAI22_X1 U1058 ( .A1(n19845), .A2(n18952), .B1(n20576), .B2(n20513), .ZN(
        n4080) );
  OAI22_X1 U1059 ( .A1(n19845), .A2(n18953), .B1(n20579), .B2(n20509), .ZN(
        n4081) );
  OAI22_X1 U1060 ( .A1(n19845), .A2(n18954), .B1(n20582), .B2(n20510), .ZN(
        n4082) );
  OAI22_X1 U1061 ( .A1(n19845), .A2(n18955), .B1(n20585), .B2(n20510), .ZN(
        n4083) );
  OAI22_X1 U1062 ( .A1(n19845), .A2(n18956), .B1(n20588), .B2(n20512), .ZN(
        n4084) );
  OAI22_X1 U1063 ( .A1(n19845), .A2(n18957), .B1(n20591), .B2(n20512), .ZN(
        n4085) );
  OAI22_X1 U1064 ( .A1(n19845), .A2(n18958), .B1(n20594), .B2(n20511), .ZN(
        n4086) );
  OAI22_X1 U1065 ( .A1(n19846), .A2(n18959), .B1(n20597), .B2(n20509), .ZN(
        n4087) );
  OAI22_X1 U1066 ( .A1(n19846), .A2(n18960), .B1(n20600), .B2(n20510), .ZN(
        n4088) );
  OAI22_X1 U1067 ( .A1(n19846), .A2(n18961), .B1(n20603), .B2(n20509), .ZN(
        n4089) );
  OAI22_X1 U1068 ( .A1(n19846), .A2(n18962), .B1(n20606), .B2(n20511), .ZN(
        n4090) );
  OAI22_X1 U1069 ( .A1(n19846), .A2(n18963), .B1(n20609), .B2(n20511), .ZN(
        n4091) );
  OAI22_X1 U1070 ( .A1(n19846), .A2(n18964), .B1(n20612), .B2(n20511), .ZN(
        n4092) );
  OAI22_X1 U1071 ( .A1(n19846), .A2(n18965), .B1(n20615), .B2(n20512), .ZN(
        n4093) );
  OAI22_X1 U1072 ( .A1(n19846), .A2(n18966), .B1(n20618), .B2(n20508), .ZN(
        n4094) );
  OAI22_X1 U1073 ( .A1(n19846), .A2(n18967), .B1(n20621), .B2(n20512), .ZN(
        n4095) );
  OAI22_X1 U1074 ( .A1(n19846), .A2(n18968), .B1(n20624), .B2(n20511), .ZN(
        n4096) );
  OAI22_X1 U1075 ( .A1(n19846), .A2(n18969), .B1(n20627), .B2(n20512), .ZN(
        n4097) );
  OAI22_X1 U1076 ( .A1(n19846), .A2(n18970), .B1(n20630), .B2(n20513), .ZN(
        n4098) );
  OAI22_X1 U1077 ( .A1(n19847), .A2(n18971), .B1(n20633), .B2(n20513), .ZN(
        n4099) );
  OAI22_X1 U1078 ( .A1(n19847), .A2(n18972), .B1(n20636), .B2(n20513), .ZN(
        n4100) );
  OAI22_X1 U1079 ( .A1(n19847), .A2(n18973), .B1(n20639), .B2(n20513), .ZN(
        n4101) );
  OAI22_X1 U1080 ( .A1(n19847), .A2(n18974), .B1(n20642), .B2(n20513), .ZN(
        n4102) );
  OAI22_X1 U1081 ( .A1(n19847), .A2(n18975), .B1(n20645), .B2(n20507), .ZN(
        n4103) );
  OAI22_X1 U1082 ( .A1(n19847), .A2(n18976), .B1(n20648), .B2(n20507), .ZN(
        n4104) );
  OAI22_X1 U1083 ( .A1(n19847), .A2(n18977), .B1(n20651), .B2(n20507), .ZN(
        n4105) );
  OAI22_X1 U1084 ( .A1(n19847), .A2(n18978), .B1(n20654), .B2(n20509), .ZN(
        n4106) );
  OAI22_X1 U1085 ( .A1(n19851), .A2(n19075), .B1(n20561), .B2(n20527), .ZN(
        n4139) );
  OAI22_X1 U1086 ( .A1(n19851), .A2(n19091), .B1(n20564), .B2(n20525), .ZN(
        n4140) );
  OAI22_X1 U1087 ( .A1(n19851), .A2(n19097), .B1(n20567), .B2(n20527), .ZN(
        n4141) );
  OAI22_X1 U1088 ( .A1(n19851), .A2(n19076), .B1(n20570), .B2(n20526), .ZN(
        n4142) );
  OAI22_X1 U1089 ( .A1(n19851), .A2(n19077), .B1(n20573), .B2(n20525), .ZN(
        n4143) );
  OAI22_X1 U1090 ( .A1(n19851), .A2(n19105), .B1(n20576), .B2(n20530), .ZN(
        n4144) );
  OAI22_X1 U1091 ( .A1(n19851), .A2(n19078), .B1(n20579), .B2(n20526), .ZN(
        n4145) );
  OAI22_X1 U1092 ( .A1(n19851), .A2(n19079), .B1(n20582), .B2(n20527), .ZN(
        n4146) );
  OAI22_X1 U1093 ( .A1(n19851), .A2(n19098), .B1(n20585), .B2(n20527), .ZN(
        n4147) );
  OAI22_X1 U1094 ( .A1(n19851), .A2(n19092), .B1(n20588), .B2(n20530), .ZN(
        n4148) );
  OAI22_X1 U1095 ( .A1(n19851), .A2(n19080), .B1(n20591), .B2(n20528), .ZN(
        n4149) );
  OAI22_X1 U1096 ( .A1(n19851), .A2(n19099), .B1(n20594), .B2(n20529), .ZN(
        n4150) );
  OAI22_X1 U1097 ( .A1(n19852), .A2(n19093), .B1(n20597), .B2(n20526), .ZN(
        n4151) );
  OAI22_X1 U1098 ( .A1(n19852), .A2(n19081), .B1(n20600), .B2(n20527), .ZN(
        n4152) );
  OAI22_X1 U1099 ( .A1(n19852), .A2(n19100), .B1(n20603), .B2(n20526), .ZN(
        n4153) );
  OAI22_X1 U1100 ( .A1(n19852), .A2(n19082), .B1(n20606), .B2(n20531), .ZN(
        n4154) );
  OAI22_X1 U1101 ( .A1(n19852), .A2(n19094), .B1(n20609), .B2(n20528), .ZN(
        n4155) );
  OAI22_X1 U1102 ( .A1(n19852), .A2(n19101), .B1(n20612), .B2(n20529), .ZN(
        n4156) );
  OAI22_X1 U1103 ( .A1(n19852), .A2(n19083), .B1(n20615), .B2(n20529), .ZN(
        n4157) );
  OAI22_X1 U1104 ( .A1(n19852), .A2(n19084), .B1(n20618), .B2(n20525), .ZN(
        n4158) );
  OAI22_X1 U1105 ( .A1(n19852), .A2(n19102), .B1(n20621), .B2(n20528), .ZN(
        n4159) );
  OAI22_X1 U1106 ( .A1(n19852), .A2(n19085), .B1(n20624), .B2(n20531), .ZN(
        n4160) );
  OAI22_X1 U1107 ( .A1(n19852), .A2(n19086), .B1(n20627), .B2(n20531), .ZN(
        n4161) );
  OAI22_X1 U1108 ( .A1(n19852), .A2(n19106), .B1(n20630), .B2(n20530), .ZN(
        n4162) );
  OAI22_X1 U1109 ( .A1(n19853), .A2(n19087), .B1(n20633), .B2(n20530), .ZN(
        n4163) );
  OAI22_X1 U1110 ( .A1(n19853), .A2(n19088), .B1(n20636), .B2(n20531), .ZN(
        n4164) );
  OAI22_X1 U1111 ( .A1(n19853), .A2(n19103), .B1(n20639), .B2(n20531), .ZN(
        n4165) );
  OAI22_X1 U1112 ( .A1(n19853), .A2(n19095), .B1(n20642), .B2(n20530), .ZN(
        n4166) );
  OAI22_X1 U1113 ( .A1(n19853), .A2(n19089), .B1(n20645), .B2(n20527), .ZN(
        n4167) );
  OAI22_X1 U1114 ( .A1(n19853), .A2(n19104), .B1(n20648), .B2(n20526), .ZN(
        n4168) );
  OAI22_X1 U1115 ( .A1(n19853), .A2(n19096), .B1(n20651), .B2(n20529), .ZN(
        n4169) );
  OAI22_X1 U1116 ( .A1(n19853), .A2(n19090), .B1(n20654), .B2(n20528), .ZN(
        n4170) );
  OAI22_X1 U1117 ( .A1(n20563), .A2(n20536), .B1(n20545), .B2(n19203), .ZN(
        n4299) );
  OAI22_X1 U1118 ( .A1(n20566), .A2(n20536), .B1(n20545), .B2(n19204), .ZN(
        n4300) );
  OAI22_X1 U1119 ( .A1(n20569), .A2(n20536), .B1(n20545), .B2(n19205), .ZN(
        n4301) );
  OAI22_X1 U1120 ( .A1(n20572), .A2(n20536), .B1(n20545), .B2(n19206), .ZN(
        n4302) );
  OAI22_X1 U1121 ( .A1(n20575), .A2(n20536), .B1(n20544), .B2(n19207), .ZN(
        n4303) );
  OAI22_X1 U1122 ( .A1(n20578), .A2(n20536), .B1(n20544), .B2(n19208), .ZN(
        n4304) );
  OAI22_X1 U1123 ( .A1(n20581), .A2(n20536), .B1(n20544), .B2(n19209), .ZN(
        n4305) );
  OAI22_X1 U1124 ( .A1(n20584), .A2(n20536), .B1(n20544), .B2(n19210), .ZN(
        n4306) );
  OAI22_X1 U1125 ( .A1(n20587), .A2(n20536), .B1(n20543), .B2(n19211), .ZN(
        n4307) );
  OAI22_X1 U1126 ( .A1(n20590), .A2(n20536), .B1(n20543), .B2(n19212), .ZN(
        n4308) );
  OAI22_X1 U1127 ( .A1(n20593), .A2(n20536), .B1(n20543), .B2(n19213), .ZN(
        n4309) );
  OAI22_X1 U1128 ( .A1(n20596), .A2(n20536), .B1(n20543), .B2(n19214), .ZN(
        n4310) );
  OAI22_X1 U1129 ( .A1(n20599), .A2(n20537), .B1(n20542), .B2(n19215), .ZN(
        n4311) );
  OAI22_X1 U1130 ( .A1(n20602), .A2(n20537), .B1(n20542), .B2(n19216), .ZN(
        n4312) );
  OAI22_X1 U1131 ( .A1(n20605), .A2(n20537), .B1(n20542), .B2(n19217), .ZN(
        n4313) );
  OAI22_X1 U1132 ( .A1(n20608), .A2(n20537), .B1(n20542), .B2(n19218), .ZN(
        n4314) );
  OAI22_X1 U1133 ( .A1(n20611), .A2(n20537), .B1(n20541), .B2(n19219), .ZN(
        n4315) );
  OAI22_X1 U1134 ( .A1(n20614), .A2(n20537), .B1(n20541), .B2(n19220), .ZN(
        n4316) );
  OAI22_X1 U1135 ( .A1(n20617), .A2(n20537), .B1(n20541), .B2(n19221), .ZN(
        n4317) );
  OAI22_X1 U1136 ( .A1(n20620), .A2(n20537), .B1(n20541), .B2(n19222), .ZN(
        n4318) );
  OAI22_X1 U1137 ( .A1(n20623), .A2(n20537), .B1(n20540), .B2(n19223), .ZN(
        n4319) );
  OAI22_X1 U1138 ( .A1(n20626), .A2(n20537), .B1(n20540), .B2(n19224), .ZN(
        n4320) );
  OAI22_X1 U1139 ( .A1(n20629), .A2(n20537), .B1(n20540), .B2(n19225), .ZN(
        n4321) );
  OAI22_X1 U1140 ( .A1(n20632), .A2(n20537), .B1(n20540), .B2(n19226), .ZN(
        n4322) );
  OAI22_X1 U1141 ( .A1(n20635), .A2(n20536), .B1(n20539), .B2(n19227), .ZN(
        n4323) );
  OAI22_X1 U1142 ( .A1(n20638), .A2(n20537), .B1(n20539), .B2(n19228), .ZN(
        n4324) );
  OAI22_X1 U1143 ( .A1(n20641), .A2(n20536), .B1(n20539), .B2(n19229), .ZN(
        n4325) );
  OAI22_X1 U1144 ( .A1(n20644), .A2(n20537), .B1(n20539), .B2(n19230), .ZN(
        n4326) );
  OAI22_X1 U1145 ( .A1(n20647), .A2(n20536), .B1(n20538), .B2(n19231), .ZN(
        n4327) );
  OAI22_X1 U1146 ( .A1(n20650), .A2(n20537), .B1(n20538), .B2(n19232), .ZN(
        n4328) );
  OAI22_X1 U1147 ( .A1(n20653), .A2(n20536), .B1(n20538), .B2(n19233), .ZN(
        n4329) );
  OAI22_X1 U1148 ( .A1(n20656), .A2(n20537), .B1(n20538), .B2(n19234), .ZN(
        n4330) );
  NAND2_X1 U1149 ( .A1(n1658), .A2(n1146), .ZN(n1657) );
  NAND2_X1 U1150 ( .A1(n1447), .A2(n1146), .ZN(n1446) );
  NAND2_X1 U1151 ( .A1(n1298), .A2(n1146), .ZN(n1297) );
  NAND2_X1 U1152 ( .A1(n1295), .A2(n1146), .ZN(n1263) );
  NAND2_X1 U1153 ( .A1(n1298), .A2(n1151), .ZN(n1335) );
  NAND2_X1 U1154 ( .A1(n1295), .A2(n1151), .ZN(n1301) );
  NAND2_X1 U1155 ( .A1(n1145), .A2(n1146), .ZN(n1079) );
  INV_X1 U1156 ( .A(ADD_RD2[0]), .ZN(n2653) );
  INV_X1 U1157 ( .A(ADD_RD1[0]), .ZN(n5707) );
  BUF_X1 U1158 ( .A(n1143), .Z(n20563) );
  BUF_X1 U1159 ( .A(n1141), .Z(n20566) );
  BUF_X1 U1160 ( .A(n1139), .Z(n20569) );
  BUF_X1 U1161 ( .A(n1137), .Z(n20572) );
  BUF_X1 U1162 ( .A(n1135), .Z(n20575) );
  BUF_X1 U1163 ( .A(n1133), .Z(n20578) );
  BUF_X1 U1164 ( .A(n1131), .Z(n20581) );
  BUF_X1 U1165 ( .A(n1129), .Z(n20584) );
  BUF_X1 U1166 ( .A(n1127), .Z(n20587) );
  BUF_X1 U1167 ( .A(n1125), .Z(n20590) );
  BUF_X1 U1168 ( .A(n1123), .Z(n20593) );
  BUF_X1 U1169 ( .A(n1121), .Z(n20596) );
  BUF_X1 U1170 ( .A(n1119), .Z(n20599) );
  BUF_X1 U1171 ( .A(n1117), .Z(n20602) );
  BUF_X1 U1172 ( .A(n1115), .Z(n20605) );
  BUF_X1 U1173 ( .A(n1113), .Z(n20608) );
  BUF_X1 U1174 ( .A(n1111), .Z(n20611) );
  BUF_X1 U1175 ( .A(n1109), .Z(n20614) );
  BUF_X1 U1176 ( .A(n1107), .Z(n20617) );
  BUF_X1 U1177 ( .A(n1105), .Z(n20620) );
  BUF_X1 U1178 ( .A(n1103), .Z(n20623) );
  BUF_X1 U1179 ( .A(n1101), .Z(n20626) );
  BUF_X1 U1180 ( .A(n1099), .Z(n20629) );
  BUF_X1 U1181 ( .A(n1097), .Z(n20632) );
  BUF_X1 U1182 ( .A(n1095), .Z(n20635) );
  BUF_X1 U1183 ( .A(n1093), .Z(n20638) );
  BUF_X1 U1184 ( .A(n1091), .Z(n20641) );
  BUF_X1 U1185 ( .A(n1089), .Z(n20644) );
  BUF_X1 U1186 ( .A(n1087), .Z(n20647) );
  BUF_X1 U1187 ( .A(n1085), .Z(n20650) );
  BUF_X1 U1188 ( .A(n1083), .Z(n20653) );
  BUF_X1 U1189 ( .A(n1080), .Z(n20656) );
  INV_X1 U1190 ( .A(ADD_RD1[4]), .ZN(n5720) );
  INV_X1 U1191 ( .A(ADD_RD2[4]), .ZN(n2690) );
  INV_X1 U1192 ( .A(ADD_RD1[3]), .ZN(n5710) );
  INV_X1 U1193 ( .A(ADD_RD2[3]), .ZN(n2675) );
  BUF_X1 U1194 ( .A(n2750), .Z(n19889) );
  INV_X1 U1195 ( .A(ADD_RD2[1]), .ZN(n2654) );
  INV_X1 U1196 ( .A(n2698), .ZN(n2694) );
  INV_X1 U1197 ( .A(n1839), .ZN(n1835) );
  INV_X1 U1198 ( .A(n5685), .ZN(n5683) );
  INV_X1 U1199 ( .A(n5640), .ZN(n5639) );
  INV_X1 U1200 ( .A(n5322), .ZN(n5321) );
  INV_X1 U1201 ( .A(n4951), .ZN(n4950) );
  INV_X1 U1202 ( .A(n4880), .ZN(n4879) );
  INV_X1 U1203 ( .A(n4762), .ZN(n4761) );
  INV_X1 U1204 ( .A(n4740), .ZN(n4739) );
  INV_X1 U1205 ( .A(n4696), .ZN(n4695) );
  INV_X1 U1206 ( .A(n4674), .ZN(n4673) );
  INV_X1 U1207 ( .A(n4630), .ZN(n4629) );
  INV_X1 U1208 ( .A(n4608), .ZN(n4607) );
  INV_X1 U1209 ( .A(n4586), .ZN(n4585) );
  INV_X1 U1210 ( .A(n4542), .ZN(n4541) );
  INV_X1 U1211 ( .A(n4520), .ZN(n4519) );
  INV_X1 U1212 ( .A(n4498), .ZN(n4497) );
  INV_X1 U1213 ( .A(n4476), .ZN(n4475) );
  INV_X1 U1214 ( .A(n2950), .ZN(n2949) );
  INV_X1 U1215 ( .A(n2928), .ZN(n2927) );
  INV_X1 U1216 ( .A(n2884), .ZN(n2883) );
  INV_X1 U1217 ( .A(n2862), .ZN(n2861) );
  INV_X1 U1218 ( .A(n2840), .ZN(n2839) );
  INV_X1 U1219 ( .A(n2796), .ZN(n2795) );
  INV_X1 U1220 ( .A(n2774), .ZN(n2773) );
  INV_X1 U1221 ( .A(n5662), .ZN(n5661) );
  INV_X1 U1222 ( .A(n4916), .ZN(n4915) );
  INV_X1 U1223 ( .A(n4718), .ZN(n4717) );
  INV_X1 U1224 ( .A(n4652), .ZN(n4651) );
  INV_X1 U1225 ( .A(n4564), .ZN(n4563) );
  INV_X1 U1226 ( .A(n2906), .ZN(n2905) );
  INV_X1 U1227 ( .A(n2818), .ZN(n2817) );
  INV_X1 U1228 ( .A(n2752), .ZN(n2751) );
  INV_X1 U1229 ( .A(n2655), .ZN(n2644) );
  INV_X1 U1230 ( .A(n2620), .ZN(n2619) );
  INV_X1 U1231 ( .A(n2595), .ZN(n2594) );
  INV_X1 U1232 ( .A(n2570), .ZN(n2569) );
  INV_X1 U1233 ( .A(n2545), .ZN(n2544) );
  INV_X1 U1234 ( .A(n2520), .ZN(n2519) );
  INV_X1 U1235 ( .A(n2495), .ZN(n2494) );
  INV_X1 U1236 ( .A(n2470), .ZN(n2469) );
  INV_X1 U1237 ( .A(n2445), .ZN(n2444) );
  INV_X1 U1238 ( .A(n2420), .ZN(n2419) );
  INV_X1 U1239 ( .A(n2395), .ZN(n2394) );
  INV_X1 U1240 ( .A(n2370), .ZN(n2369) );
  INV_X1 U1241 ( .A(n2345), .ZN(n2344) );
  INV_X1 U1242 ( .A(n2320), .ZN(n2319) );
  INV_X1 U1243 ( .A(n2295), .ZN(n2294) );
  INV_X1 U1244 ( .A(n2270), .ZN(n2269) );
  INV_X1 U1245 ( .A(n2245), .ZN(n2244) );
  INV_X1 U1246 ( .A(n2220), .ZN(n2219) );
  INV_X1 U1247 ( .A(n2195), .ZN(n2194) );
  INV_X1 U1248 ( .A(n2170), .ZN(n2169) );
  INV_X1 U1249 ( .A(n2145), .ZN(n2144) );
  INV_X1 U1250 ( .A(n2120), .ZN(n2119) );
  INV_X1 U1251 ( .A(n2095), .ZN(n2094) );
  INV_X1 U1252 ( .A(n2070), .ZN(n2069) );
  INV_X1 U1253 ( .A(n2045), .ZN(n2044) );
  INV_X1 U1254 ( .A(n2020), .ZN(n2019) );
  INV_X1 U1255 ( .A(n1995), .ZN(n1994) );
  INV_X1 U1256 ( .A(n1970), .ZN(n1969) );
  INV_X1 U1257 ( .A(n1945), .ZN(n1944) );
  INV_X1 U1258 ( .A(n1920), .ZN(n1919) );
  INV_X1 U1259 ( .A(n1895), .ZN(n1894) );
  INV_X1 U1260 ( .A(ADD_RD1[1]), .ZN(n5718) );
  INV_X1 U1261 ( .A(ADD_RD2[2]), .ZN(n2689) );
  OAI22_X1 U1262 ( .A1(n19259), .A2(n19949), .B1(n18907), .B2(n19958), .ZN(
        n4495) );
  OAI22_X1 U1263 ( .A1(n19260), .A2(n19949), .B1(n18908), .B2(n19958), .ZN(
        n4473) );
  OAI22_X1 U1264 ( .A1(n19261), .A2(n19951), .B1(n18909), .B2(n19959), .ZN(
        n2947) );
  OAI22_X1 U1265 ( .A1(n19262), .A2(n19951), .B1(n18911), .B2(n19957), .ZN(
        n2903) );
  OAI22_X1 U1266 ( .A1(n19263), .A2(n19951), .B1(n18912), .B2(n19956), .ZN(
        n2881) );
  OAI22_X1 U1267 ( .A1(n19264), .A2(n19950), .B1(n18913), .B2(n19959), .ZN(
        n2859) );
  OAI22_X1 U1268 ( .A1(n19265), .A2(n19951), .B1(n18910), .B2(n19959), .ZN(
        n2925) );
  OAI22_X1 U1269 ( .A1(n19266), .A2(n19949), .B1(n18914), .B2(n19957), .ZN(
        n2837) );
  OAI22_X1 U1270 ( .A1(n18875), .A2(n19919), .B1(n19127), .B2(n19927), .ZN(
        n4496) );
  OAI22_X1 U1271 ( .A1(n18876), .A2(n19919), .B1(n19128), .B2(n19927), .ZN(
        n4474) );
  OAI22_X1 U1272 ( .A1(n18877), .A2(n19919), .B1(n19129), .B2(n19926), .ZN(
        n2948) );
  OAI22_X1 U1273 ( .A1(n18878), .A2(n19919), .B1(n19131), .B2(n19925), .ZN(
        n2904) );
  OAI22_X1 U1274 ( .A1(n18879), .A2(n19919), .B1(n19132), .B2(n19927), .ZN(
        n2882) );
  OAI22_X1 U1275 ( .A1(n18880), .A2(n19917), .B1(n19133), .B2(n19927), .ZN(
        n2860) );
  OAI22_X1 U1276 ( .A1(n18881), .A2(n19918), .B1(n19130), .B2(n19927), .ZN(
        n2926) );
  OAI22_X1 U1277 ( .A1(n18882), .A2(n19917), .B1(n19134), .B2(n19926), .ZN(
        n2838) );
  BUF_X1 U1278 ( .A(n1078), .Z(n20668) );
  BUF_X1 U1279 ( .A(n1078), .Z(n20667) );
  BUF_X1 U1280 ( .A(n1078), .Z(n20666) );
  NAND2_X1 U1281 ( .A1(n1225), .A2(n1145), .ZN(n20533) );
  NAND2_X1 U1282 ( .A1(n1225), .A2(n1145), .ZN(n1226) );
  NAND2_X1 U1283 ( .A1(n1188), .A2(n1145), .ZN(n20535) );
  NAND2_X1 U1284 ( .A1(n1188), .A2(n1145), .ZN(n1190) );
  NAND2_X1 U1285 ( .A1(n1658), .A2(n1225), .ZN(n1833) );
  NAND2_X1 U1286 ( .A1(n1655), .A2(n1225), .ZN(n1799) );
  NAND2_X1 U1287 ( .A1(n1658), .A2(n1188), .ZN(n1764) );
  NAND2_X1 U1288 ( .A1(n1655), .A2(n1188), .ZN(n1730) );
  NAND2_X1 U1289 ( .A1(n1447), .A2(n1225), .ZN(n1589) );
  NAND2_X1 U1290 ( .A1(n1447), .A2(n1188), .ZN(n1520) );
  NAND2_X1 U1291 ( .A1(n1444), .A2(n1188), .ZN(n1517) );
  NAND2_X1 U1292 ( .A1(n1295), .A2(n1225), .ZN(n20473) );
  NAND2_X1 U1293 ( .A1(n1295), .A2(n1225), .ZN(n1405) );
  NAND2_X1 U1294 ( .A1(n1295), .A2(n1188), .ZN(n20489) );
  NAND2_X1 U1295 ( .A1(n1295), .A2(n1188), .ZN(n1368) );
  NAND2_X1 U1296 ( .A1(n1655), .A2(n1146), .ZN(n1623) );
  NAND2_X1 U1297 ( .A1(n1444), .A2(n1146), .ZN(n1443) );
  NAND2_X1 U1298 ( .A1(n1658), .A2(n1151), .ZN(n1695) );
  NAND2_X1 U1299 ( .A1(n1655), .A2(n1151), .ZN(n1661) );
  NAND2_X1 U1300 ( .A1(n1447), .A2(n1151), .ZN(n1484) );
  NAND2_X1 U1301 ( .A1(n1444), .A2(n1151), .ZN(n1450) );
  BUF_X1 U1302 ( .A(n19882), .Z(n19884) );
  BUF_X1 U1303 ( .A(n19882), .Z(n19885) );
  BUF_X1 U1304 ( .A(n19883), .Z(n19886) );
  AND2_X1 U1305 ( .A1(n1586), .A2(n1150), .ZN(n1444) );
  BUF_X1 U1306 ( .A(n19883), .Z(n19887) );
  BUF_X1 U1307 ( .A(n2750), .Z(n19888) );
  BUF_X1 U1308 ( .A(n20757), .Z(n20686) );
  BUF_X1 U1309 ( .A(n20758), .Z(n20757) );
  BUF_X1 U1310 ( .A(n19875), .Z(n19878) );
  BUF_X1 U1311 ( .A(n19874), .Z(n19876) );
  BUF_X1 U1312 ( .A(n19874), .Z(n19877) );
  BUF_X1 U1313 ( .A(n19866), .Z(n19868) );
  BUF_X1 U1314 ( .A(n19866), .Z(n19869) );
  BUF_X1 U1315 ( .A(n19867), .Z(n19870) );
  BUF_X1 U1316 ( .A(n2697), .Z(n19880) );
  BUF_X1 U1317 ( .A(n19875), .Z(n19879) );
  BUF_X1 U1318 ( .A(n19867), .Z(n19871) );
  BUF_X1 U1319 ( .A(n1838), .Z(n19872) );
  BUF_X1 U1320 ( .A(n2697), .Z(n19881) );
  BUF_X1 U1321 ( .A(n1838), .Z(n19873) );
  NAND2_X1 U1322 ( .A1(n19881), .A2(n5685), .ZN(n3086) );
  NAND2_X1 U1323 ( .A1(n19878), .A2(n5640), .ZN(n3098) );
  NAND2_X1 U1324 ( .A1(n19879), .A2(n5322), .ZN(n3104) );
  NAND2_X1 U1325 ( .A1(n19880), .A2(n4951), .ZN(n3110) );
  NAND2_X1 U1326 ( .A1(n19877), .A2(n4880), .ZN(n3122) );
  NAND2_X1 U1327 ( .A1(n19878), .A2(n4762), .ZN(n3128) );
  NAND2_X1 U1328 ( .A1(n19881), .A2(n4740), .ZN(n3134) );
  NAND2_X1 U1329 ( .A1(n19877), .A2(n4696), .ZN(n3146) );
  NAND2_X1 U1330 ( .A1(n19880), .A2(n4674), .ZN(n3152) );
  NAND2_X1 U1331 ( .A1(n19880), .A2(n4630), .ZN(n3164) );
  NAND2_X1 U1332 ( .A1(n19878), .A2(n4608), .ZN(n3170) );
  NAND2_X1 U1333 ( .A1(n19879), .A2(n4586), .ZN(n3176) );
  NAND2_X1 U1334 ( .A1(n19881), .A2(n4542), .ZN(n3188) );
  NAND2_X1 U1335 ( .A1(n19881), .A2(n4520), .ZN(n3194) );
  NAND2_X1 U1336 ( .A1(n19876), .A2(n4498), .ZN(n3200) );
  NAND2_X1 U1337 ( .A1(n19881), .A2(n4476), .ZN(n3206) );
  NAND2_X1 U1338 ( .A1(n19876), .A2(n2950), .ZN(n3212) );
  NAND2_X1 U1339 ( .A1(n19877), .A2(n2928), .ZN(n3218) );
  NAND2_X1 U1340 ( .A1(n19877), .A2(n2884), .ZN(n3230) );
  NAND2_X1 U1341 ( .A1(n19878), .A2(n2862), .ZN(n3236) );
  NAND2_X1 U1342 ( .A1(n19878), .A2(n2840), .ZN(n3242) );
  NAND2_X1 U1343 ( .A1(n19880), .A2(n2796), .ZN(n3254) );
  NAND2_X1 U1344 ( .A1(n19877), .A2(n2774), .ZN(n3260) );
  NAND2_X1 U1345 ( .A1(n19880), .A2(n2698), .ZN(n3272) );
  NAND2_X1 U1346 ( .A1(n19876), .A2(n5662), .ZN(n3092) );
  NAND2_X1 U1347 ( .A1(n19879), .A2(n4916), .ZN(n3116) );
  NAND2_X1 U1348 ( .A1(n19876), .A2(n4718), .ZN(n3140) );
  NAND2_X1 U1349 ( .A1(n19879), .A2(n4652), .ZN(n3158) );
  NAND2_X1 U1350 ( .A1(n19880), .A2(n4564), .ZN(n3182) );
  NAND2_X1 U1351 ( .A1(n19876), .A2(n2906), .ZN(n3224) );
  NAND2_X1 U1352 ( .A1(n19879), .A2(n2818), .ZN(n3248) );
  NAND2_X1 U1353 ( .A1(n19879), .A2(n2752), .ZN(n3266) );
  NAND2_X1 U1354 ( .A1(n19873), .A2(n2655), .ZN(n3276) );
  NAND2_X1 U1355 ( .A1(n19868), .A2(n2620), .ZN(n3281) );
  NAND2_X1 U1356 ( .A1(n19870), .A2(n2595), .ZN(n3286) );
  NAND2_X1 U1357 ( .A1(n19871), .A2(n2570), .ZN(n3291) );
  NAND2_X1 U1358 ( .A1(n19872), .A2(n2545), .ZN(n3296) );
  NAND2_X1 U1359 ( .A1(n19871), .A2(n2520), .ZN(n3301) );
  NAND2_X1 U1360 ( .A1(n19869), .A2(n2495), .ZN(n3306) );
  NAND2_X1 U1361 ( .A1(n19870), .A2(n2470), .ZN(n3311) );
  NAND2_X1 U1362 ( .A1(n19873), .A2(n2445), .ZN(n3316) );
  NAND2_X1 U1363 ( .A1(n19868), .A2(n2420), .ZN(n3321) );
  NAND2_X1 U1364 ( .A1(n19869), .A2(n2395), .ZN(n3326) );
  NAND2_X1 U1365 ( .A1(n19872), .A2(n2370), .ZN(n3331) );
  NAND2_X1 U1366 ( .A1(n19871), .A2(n2345), .ZN(n3336) );
  NAND2_X1 U1367 ( .A1(n19872), .A2(n2320), .ZN(n3341) );
  NAND2_X1 U1368 ( .A1(n19870), .A2(n2295), .ZN(n3346) );
  NAND2_X1 U1369 ( .A1(n19871), .A2(n2270), .ZN(n3351) );
  NAND2_X1 U1370 ( .A1(n19872), .A2(n2245), .ZN(n3356) );
  NAND2_X1 U1371 ( .A1(n19873), .A2(n2220), .ZN(n3361) );
  NAND2_X1 U1372 ( .A1(n19873), .A2(n2195), .ZN(n3366) );
  NAND2_X1 U1373 ( .A1(n19868), .A2(n2170), .ZN(n3371) );
  NAND2_X1 U1374 ( .A1(n19873), .A2(n2145), .ZN(n3376) );
  NAND2_X1 U1375 ( .A1(n19868), .A2(n2120), .ZN(n3381) );
  NAND2_X1 U1376 ( .A1(n19869), .A2(n2095), .ZN(n3386) );
  NAND2_X1 U1377 ( .A1(n19868), .A2(n2070), .ZN(n3391) );
  NAND2_X1 U1378 ( .A1(n19869), .A2(n2045), .ZN(n3396) );
  NAND2_X1 U1379 ( .A1(n19870), .A2(n2020), .ZN(n3401) );
  NAND2_X1 U1380 ( .A1(n19870), .A2(n1995), .ZN(n3406) );
  NAND2_X1 U1381 ( .A1(n19871), .A2(n1970), .ZN(n3411) );
  NAND2_X1 U1382 ( .A1(n19872), .A2(n1945), .ZN(n3416) );
  NAND2_X1 U1383 ( .A1(n19869), .A2(n1920), .ZN(n3421) );
  NAND2_X1 U1384 ( .A1(n19871), .A2(n1895), .ZN(n3426) );
  NAND2_X1 U1385 ( .A1(n19872), .A2(n1839), .ZN(n3431) );
  BUF_X1 U1386 ( .A(n20758), .Z(n20752) );
  BUF_X1 U1387 ( .A(n20758), .Z(n20750) );
  BUF_X1 U1388 ( .A(n20758), .Z(n20747) );
  BUF_X1 U1389 ( .A(n20758), .Z(n20754) );
  BUF_X1 U1390 ( .A(n20758), .Z(n20756) );
  BUF_X1 U1391 ( .A(n20758), .Z(n20753) );
  BUF_X1 U1392 ( .A(n20758), .Z(n20748) );
  BUF_X1 U1393 ( .A(n20758), .Z(n20755) );
  BUF_X1 U1394 ( .A(n20758), .Z(n20751) );
  BUF_X1 U1395 ( .A(n20758), .Z(n20749) );
  INV_X1 U1396 ( .A(DATAIN[0]), .ZN(n1143) );
  INV_X1 U1397 ( .A(DATAIN[1]), .ZN(n1141) );
  INV_X1 U1398 ( .A(DATAIN[2]), .ZN(n1139) );
  INV_X1 U1399 ( .A(DATAIN[3]), .ZN(n1137) );
  INV_X1 U1400 ( .A(DATAIN[4]), .ZN(n1135) );
  INV_X1 U1401 ( .A(DATAIN[5]), .ZN(n1133) );
  INV_X1 U1402 ( .A(DATAIN[6]), .ZN(n1131) );
  INV_X1 U1403 ( .A(DATAIN[7]), .ZN(n1129) );
  INV_X1 U1404 ( .A(DATAIN[8]), .ZN(n1127) );
  INV_X1 U1405 ( .A(DATAIN[9]), .ZN(n1125) );
  INV_X1 U1406 ( .A(DATAIN[10]), .ZN(n1123) );
  INV_X1 U1407 ( .A(DATAIN[11]), .ZN(n1121) );
  INV_X1 U1408 ( .A(DATAIN[12]), .ZN(n1119) );
  INV_X1 U1409 ( .A(DATAIN[13]), .ZN(n1117) );
  INV_X1 U1410 ( .A(DATAIN[14]), .ZN(n1115) );
  INV_X1 U1411 ( .A(DATAIN[15]), .ZN(n1113) );
  INV_X1 U1412 ( .A(DATAIN[16]), .ZN(n1111) );
  INV_X1 U1413 ( .A(DATAIN[17]), .ZN(n1109) );
  INV_X1 U1414 ( .A(DATAIN[18]), .ZN(n1107) );
  INV_X1 U1415 ( .A(DATAIN[19]), .ZN(n1105) );
  INV_X1 U1416 ( .A(DATAIN[20]), .ZN(n1103) );
  INV_X1 U1417 ( .A(DATAIN[21]), .ZN(n1101) );
  INV_X1 U1418 ( .A(DATAIN[22]), .ZN(n1099) );
  INV_X1 U1419 ( .A(DATAIN[23]), .ZN(n1097) );
  INV_X1 U1420 ( .A(DATAIN[24]), .ZN(n1095) );
  INV_X1 U1421 ( .A(DATAIN[25]), .ZN(n1093) );
  INV_X1 U1422 ( .A(DATAIN[26]), .ZN(n1091) );
  INV_X1 U1423 ( .A(DATAIN[27]), .ZN(n1089) );
  INV_X1 U1424 ( .A(DATAIN[28]), .ZN(n1087) );
  INV_X1 U1425 ( .A(DATAIN[29]), .ZN(n1085) );
  INV_X1 U1426 ( .A(DATAIN[30]), .ZN(n1083) );
  INV_X1 U1427 ( .A(DATAIN[31]), .ZN(n1080) );
  NOR4_X1 U1428 ( .A1(n2660), .A2(n2661), .A3(n2662), .A4(n2663), .ZN(n2659)
         );
  OAI221_X1 U1429 ( .B1(n8657), .B2(n20233), .C1(n19395), .C2(n20236), .A(
        n2678), .ZN(n2660) );
  OAI221_X1 U1430 ( .B1(n19075), .B2(n20285), .C1(n8454), .C2(n20288), .A(
        n2670), .ZN(n2662) );
  OAI221_X1 U1431 ( .B1(n19299), .B2(n20299), .C1(n5541), .C2(n20307), .A(
        n2664), .ZN(n2663) );
  NOR4_X1 U1432 ( .A1(n2625), .A2(n2626), .A3(n2627), .A4(n2628), .ZN(n2624)
         );
  OAI221_X1 U1433 ( .B1(n8658), .B2(n20233), .C1(n19396), .C2(n20236), .A(
        n2634), .ZN(n2625) );
  OAI221_X1 U1434 ( .B1(n19091), .B2(n20286), .C1(n8455), .C2(n20289), .A(
        n2630), .ZN(n2627) );
  OAI221_X1 U1435 ( .B1(n19300), .B2(n20300), .C1(n5542), .C2(n20308), .A(
        n2629), .ZN(n2628) );
  NOR4_X1 U1436 ( .A1(n2575), .A2(n2576), .A3(n2577), .A4(n2578), .ZN(n2574)
         );
  OAI221_X1 U1437 ( .B1(n8660), .B2(n20233), .C1(n19397), .C2(n20236), .A(
        n2584), .ZN(n2575) );
  OAI221_X1 U1438 ( .B1(n19076), .B2(n20285), .C1(n8456), .C2(n20289), .A(
        n2580), .ZN(n2577) );
  OAI221_X1 U1439 ( .B1(n19301), .B2(n20300), .C1(n5544), .C2(n20308), .A(
        n2579), .ZN(n2578) );
  NOR4_X1 U1440 ( .A1(n2550), .A2(n2551), .A3(n2552), .A4(n2553), .ZN(n2549)
         );
  OAI221_X1 U1441 ( .B1(n8661), .B2(n20229), .C1(n19398), .C2(n20237), .A(
        n2559), .ZN(n2550) );
  OAI221_X1 U1442 ( .B1(n19077), .B2(n20286), .C1(n8457), .C2(n20290), .A(
        n2555), .ZN(n2552) );
  OAI221_X1 U1443 ( .B1(n19302), .B2(n20300), .C1(n5545), .C2(n20309), .A(
        n2554), .ZN(n2553) );
  NOR4_X1 U1444 ( .A1(n2500), .A2(n2501), .A3(n2502), .A4(n2503), .ZN(n2499)
         );
  OAI221_X1 U1445 ( .B1(n8663), .B2(n20232), .C1(n19399), .C2(n20240), .A(
        n2509), .ZN(n2500) );
  OAI221_X1 U1446 ( .B1(n19078), .B2(n20285), .C1(n8461), .C2(n20290), .A(
        n2505), .ZN(n2502) );
  OAI221_X1 U1447 ( .B1(n19303), .B2(n20303), .C1(n5547), .C2(n20309), .A(
        n2504), .ZN(n2503) );
  NOR4_X1 U1448 ( .A1(n2475), .A2(n2476), .A3(n2477), .A4(n2478), .ZN(n2474)
         );
  OAI221_X1 U1449 ( .B1(n8664), .B2(n20229), .C1(n19400), .C2(n20238), .A(
        n2484), .ZN(n2475) );
  OAI221_X1 U1450 ( .B1(n19079), .B2(n20286), .C1(n8462), .C2(n20291), .A(
        n2480), .ZN(n2477) );
  OAI221_X1 U1451 ( .B1(n19304), .B2(n20301), .C1(n5548), .C2(n20310), .A(
        n2479), .ZN(n2478) );
  NOR4_X1 U1452 ( .A1(n2425), .A2(n2426), .A3(n2427), .A4(n2428), .ZN(n2424)
         );
  OAI221_X1 U1453 ( .B1(n8665), .B2(n20234), .C1(n19401), .C2(n20236), .A(
        n2434), .ZN(n2425) );
  OAI221_X1 U1454 ( .B1(n19092), .B2(n20285), .C1(n8463), .C2(n20293), .A(
        n2430), .ZN(n2427) );
  OAI221_X1 U1455 ( .B1(n19305), .B2(n20300), .C1(n5550), .C2(n20312), .A(
        n2429), .ZN(n2428) );
  NOR4_X1 U1456 ( .A1(n2400), .A2(n2401), .A3(n2402), .A4(n2403), .ZN(n2399)
         );
  OAI221_X1 U1457 ( .B1(n8666), .B2(n20230), .C1(n19402), .C2(n20239), .A(
        n2409), .ZN(n2400) );
  OAI221_X1 U1458 ( .B1(n19080), .B2(n20286), .C1(n8464), .C2(n20288), .A(
        n2405), .ZN(n2402) );
  OAI221_X1 U1459 ( .B1(n19306), .B2(n20302), .C1(n5551), .C2(n20307), .A(
        n2404), .ZN(n2403) );
  NOR4_X1 U1460 ( .A1(n2350), .A2(n2351), .A3(n2352), .A4(n2353), .ZN(n2349)
         );
  OAI221_X1 U1461 ( .B1(n8673), .B2(n20228), .C1(n19403), .C2(n20237), .A(
        n2359), .ZN(n2350) );
  OAI221_X1 U1462 ( .B1(n19093), .B2(n20285), .C1(n8465), .C2(n20292), .A(
        n2355), .ZN(n2352) );
  OAI221_X1 U1463 ( .B1(n19307), .B2(n20300), .C1(n5553), .C2(n20311), .A(
        n2354), .ZN(n2353) );
  NOR4_X1 U1464 ( .A1(n2325), .A2(n2326), .A3(n2327), .A4(n2328), .ZN(n2324)
         );
  OAI221_X1 U1465 ( .B1(n8674), .B2(n20228), .C1(n19404), .C2(n20238), .A(
        n2334), .ZN(n2325) );
  OAI221_X1 U1466 ( .B1(n19081), .B2(n20286), .C1(n8466), .C2(n20293), .A(
        n2330), .ZN(n2327) );
  OAI221_X1 U1467 ( .B1(n19308), .B2(n20299), .C1(n5554), .C2(n20312), .A(
        n2329), .ZN(n2328) );
  NOR4_X1 U1468 ( .A1(n2275), .A2(n2276), .A3(n2277), .A4(n2278), .ZN(n2274)
         );
  OAI221_X1 U1469 ( .B1(n8667), .B2(n20229), .C1(n19405), .C2(n20238), .A(
        n2284), .ZN(n2275) );
  OAI221_X1 U1470 ( .B1(n19082), .B2(n20285), .C1(n8470), .C2(n20291), .A(
        n2280), .ZN(n2277) );
  OAI221_X1 U1471 ( .B1(n19309), .B2(n20301), .C1(n5556), .C2(n20310), .A(
        n2279), .ZN(n2278) );
  NOR4_X1 U1472 ( .A1(n2250), .A2(n2251), .A3(n2252), .A4(n2253), .ZN(n2249)
         );
  OAI221_X1 U1473 ( .B1(n8668), .B2(n20230), .C1(n19406), .C2(n20242), .A(
        n2259), .ZN(n2250) );
  OAI221_X1 U1474 ( .B1(n19094), .B2(n20286), .C1(n8471), .C2(n20292), .A(
        n2255), .ZN(n2252) );
  OAI221_X1 U1475 ( .B1(n19310), .B2(n20305), .C1(n5557), .C2(n20311), .A(
        n2254), .ZN(n2253) );
  NOR4_X1 U1476 ( .A1(n2200), .A2(n2201), .A3(n2202), .A4(n2203), .ZN(n2199)
         );
  OAI221_X1 U1477 ( .B1(n8669), .B2(n20230), .C1(n19407), .C2(n20239), .A(
        n2209), .ZN(n2200) );
  OAI221_X1 U1478 ( .B1(n19083), .B2(n20285), .C1(n8472), .C2(n20288), .A(
        n2205), .ZN(n2202) );
  OAI221_X1 U1479 ( .B1(n19311), .B2(n20302), .C1(n5559), .C2(n20307), .A(
        n2204), .ZN(n2203) );
  NOR4_X1 U1480 ( .A1(n2175), .A2(n2176), .A3(n2177), .A4(n2178), .ZN(n2174)
         );
  OAI221_X1 U1481 ( .B1(n8670), .B2(n20231), .C1(n19408), .C2(n20240), .A(
        n2184), .ZN(n2175) );
  OAI221_X1 U1482 ( .B1(n19084), .B2(n20286), .C1(n8458), .C2(n20289), .A(
        n2180), .ZN(n2177) );
  OAI221_X1 U1483 ( .B1(n19312), .B2(n20303), .C1(n5560), .C2(n20308), .A(
        n2179), .ZN(n2178) );
  NOR4_X1 U1484 ( .A1(n2125), .A2(n2126), .A3(n2127), .A4(n2128), .ZN(n2124)
         );
  OAI221_X1 U1485 ( .B1(n8678), .B2(n20232), .C1(n19409), .C2(n20240), .A(
        n2134), .ZN(n2125) );
  OAI221_X1 U1486 ( .B1(n19313), .B2(n20303), .C1(n5562), .C2(n20308), .A(
        n2129), .ZN(n2128) );
  OAI221_X1 U1487 ( .B1(n19085), .B2(n20285), .C1(n8475), .C2(n20289), .A(
        n2130), .ZN(n2127) );
  NOR4_X1 U1488 ( .A1(n2100), .A2(n2101), .A3(n2102), .A4(n2103), .ZN(n2099)
         );
  OAI221_X1 U1489 ( .B1(n8679), .B2(n20232), .C1(n19410), .C2(n20241), .A(
        n2109), .ZN(n2100) );
  OAI221_X1 U1490 ( .B1(n19314), .B2(n20304), .C1(n5563), .C2(n20309), .A(
        n2104), .ZN(n2103) );
  OAI221_X1 U1491 ( .B1(n19086), .B2(n20286), .C1(n8476), .C2(n20290), .A(
        n2105), .ZN(n2102) );
  NOR4_X1 U1492 ( .A1(n2050), .A2(n2051), .A3(n2052), .A4(n2053), .ZN(n2049)
         );
  OAI221_X1 U1493 ( .B1(n8681), .B2(n20233), .C1(n19411), .C2(n20242), .A(
        n2059), .ZN(n2050) );
  OAI221_X1 U1494 ( .B1(n19315), .B2(n20305), .C1(n5564), .C2(n20309), .A(
        n2054), .ZN(n2053) );
  OAI221_X1 U1495 ( .B1(n19087), .B2(n20285), .C1(n8478), .C2(n20290), .A(
        n2055), .ZN(n2052) );
  NOR4_X1 U1496 ( .A1(n2025), .A2(n2026), .A3(n2027), .A4(n2028), .ZN(n2024)
         );
  OAI221_X1 U1497 ( .B1(n8682), .B2(n20234), .C1(n19412), .C2(n20242), .A(
        n2034), .ZN(n2025) );
  OAI221_X1 U1498 ( .B1(n19316), .B2(n20305), .C1(n5565), .C2(n20310), .A(
        n2029), .ZN(n2028) );
  OAI221_X1 U1499 ( .B1(n19088), .B2(n20286), .C1(n8479), .C2(n20291), .A(
        n2030), .ZN(n2027) );
  NOR4_X1 U1500 ( .A1(n1975), .A2(n1976), .A3(n1977), .A4(n1978), .ZN(n1974)
         );
  OAI221_X1 U1501 ( .B1(n8683), .B2(n20234), .C1(n19413), .C2(n20242), .A(
        n1984), .ZN(n1975) );
  OAI221_X1 U1502 ( .B1(n19317), .B2(n20305), .C1(n5567), .C2(n20312), .A(
        n1979), .ZN(n1978) );
  OAI221_X1 U1503 ( .B1(n19095), .B2(n20285), .C1(n8480), .C2(n20293), .A(
        n1980), .ZN(n1977) );
  NOR4_X1 U1504 ( .A1(n1950), .A2(n1951), .A3(n1952), .A4(n1953), .ZN(n1949)
         );
  OAI221_X1 U1505 ( .B1(n8684), .B2(n20233), .C1(n19414), .C2(n20236), .A(
        n1959), .ZN(n1950) );
  OAI221_X1 U1506 ( .B1(n19089), .B2(n20286), .C1(n8481), .C2(n20288), .A(
        n1955), .ZN(n1952) );
  OAI221_X1 U1507 ( .B1(n19318), .B2(n20299), .C1(n5568), .C2(n20307), .A(
        n1954), .ZN(n1953) );
  NOR4_X1 U1508 ( .A1(n1900), .A2(n1901), .A3(n1902), .A4(n1903), .ZN(n1899)
         );
  OAI221_X1 U1509 ( .B1(n8688), .B2(n20229), .C1(n19415), .C2(n20237), .A(
        n1909), .ZN(n1900) );
  OAI221_X1 U1510 ( .B1(n19096), .B2(n20285), .C1(n8484), .C2(n20292), .A(
        n1905), .ZN(n1902) );
  OAI221_X1 U1511 ( .B1(n19319), .B2(n20301), .C1(n5570), .C2(n20311), .A(
        n1904), .ZN(n1903) );
  NOR4_X1 U1512 ( .A1(n1844), .A2(n1845), .A3(n1846), .A4(n1847), .ZN(n1843)
         );
  OAI221_X1 U1513 ( .B1(n8685), .B2(n20234), .C1(n19416), .C2(n20242), .A(
        n1867), .ZN(n1844) );
  OAI221_X1 U1514 ( .B1(n19090), .B2(n20286), .C1(n8485), .C2(n20293), .A(
        n1855), .ZN(n1846) );
  OAI221_X1 U1515 ( .B1(n19320), .B2(n20305), .C1(n5571), .C2(n20312), .A(
        n1850), .ZN(n1847) );
  NOR4_X1 U1516 ( .A1(n2600), .A2(n2601), .A3(n2602), .A4(n2603), .ZN(n2599)
         );
  OAI221_X1 U1517 ( .B1(n8659), .B2(n20228), .C1(n19417), .C2(n20237), .A(
        n2609), .ZN(n2600) );
  OAI221_X1 U1518 ( .B1(n19097), .B2(n1853), .C1(n8459), .C2(n20288), .A(n2605), .ZN(n2602) );
  OAI221_X1 U1519 ( .B1(n19321), .B2(n20299), .C1(n5543), .C2(n20307), .A(
        n2604), .ZN(n2603) );
  NOR4_X1 U1520 ( .A1(n2525), .A2(n2526), .A3(n2527), .A4(n2528), .ZN(n2524)
         );
  OAI221_X1 U1521 ( .B1(n8662), .B2(n20228), .C1(n19418), .C2(n20238), .A(
        n2534), .ZN(n2525) );
  OAI221_X1 U1522 ( .B1(n19105), .B2(n1853), .C1(n8460), .C2(n20291), .A(n2530), .ZN(n2527) );
  OAI221_X1 U1523 ( .B1(n19322), .B2(n20301), .C1(n5546), .C2(n20310), .A(
        n2529), .ZN(n2528) );
  NOR4_X1 U1524 ( .A1(n2450), .A2(n2451), .A3(n2452), .A4(n2453), .ZN(n2449)
         );
  OAI221_X1 U1525 ( .B1(n8671), .B2(n20231), .C1(n19419), .C2(n20237), .A(
        n2459), .ZN(n2450) );
  OAI221_X1 U1526 ( .B1(n19098), .B2(n1853), .C1(n8467), .C2(n20292), .A(n2455), .ZN(n2452) );
  OAI221_X1 U1527 ( .B1(n19323), .B2(n20299), .C1(n5549), .C2(n20311), .A(
        n2454), .ZN(n2453) );
  NOR4_X1 U1528 ( .A1(n2375), .A2(n2376), .A3(n2377), .A4(n2378), .ZN(n2374)
         );
  OAI221_X1 U1529 ( .B1(n8672), .B2(n20231), .C1(n19420), .C2(n20240), .A(
        n2384), .ZN(n2375) );
  OAI221_X1 U1530 ( .B1(n19099), .B2(n1853), .C1(n8468), .C2(n20289), .A(n2380), .ZN(n2377) );
  OAI221_X1 U1531 ( .B1(n19324), .B2(n20303), .C1(n5552), .C2(n20308), .A(
        n2379), .ZN(n2378) );
  NOR4_X1 U1532 ( .A1(n2300), .A2(n2301), .A3(n2302), .A4(n2303), .ZN(n2299)
         );
  OAI221_X1 U1533 ( .B1(n8675), .B2(n20229), .C1(n19421), .C2(n20241), .A(
        n2309), .ZN(n2300) );
  OAI221_X1 U1534 ( .B1(n19100), .B2(n1853), .C1(n8469), .C2(n20290), .A(n2305), .ZN(n2302) );
  OAI221_X1 U1535 ( .B1(n19325), .B2(n20302), .C1(n5555), .C2(n20309), .A(
        n2304), .ZN(n2303) );
  NOR4_X1 U1536 ( .A1(n2225), .A2(n2226), .A3(n2227), .A4(n2228), .ZN(n2224)
         );
  OAI221_X1 U1537 ( .B1(n8676), .B2(n20233), .C1(n19422), .C2(n20239), .A(
        n2234), .ZN(n2225) );
  OAI221_X1 U1538 ( .B1(n19101), .B2(n1853), .C1(n8473), .C2(n20293), .A(n2230), .ZN(n2227) );
  OAI221_X1 U1539 ( .B1(n19326), .B2(n20304), .C1(n5558), .C2(n20312), .A(
        n2229), .ZN(n2228) );
  NOR4_X1 U1540 ( .A1(n2150), .A2(n2151), .A3(n2152), .A4(n2153), .ZN(n2149)
         );
  OAI221_X1 U1541 ( .B1(n8677), .B2(n20231), .C1(n19423), .C2(n20241), .A(
        n2159), .ZN(n2150) );
  OAI221_X1 U1542 ( .B1(n19327), .B2(n20304), .C1(n5561), .C2(n20307), .A(
        n2154), .ZN(n2153) );
  OAI221_X1 U1543 ( .B1(n19102), .B2(n1853), .C1(n8474), .C2(n20288), .A(n2155), .ZN(n2152) );
  NOR4_X1 U1544 ( .A1(n2075), .A2(n2076), .A3(n2077), .A4(n2078), .ZN(n2074)
         );
  OAI221_X1 U1545 ( .B1(n8680), .B2(n20232), .C1(n19424), .C2(n20239), .A(
        n2084), .ZN(n2075) );
  OAI221_X1 U1546 ( .B1(n19328), .B2(n20302), .C1(n5477), .C2(n20310), .A(
        n2079), .ZN(n2078) );
  OAI221_X1 U1547 ( .B1(n19106), .B2(n1853), .C1(n8477), .C2(n20291), .A(n2080), .ZN(n2077) );
  NOR4_X1 U1548 ( .A1(n2000), .A2(n2001), .A3(n2002), .A4(n2003), .ZN(n1999)
         );
  OAI221_X1 U1549 ( .B1(n8686), .B2(n20230), .C1(n19425), .C2(n20241), .A(
        n2009), .ZN(n2000) );
  OAI221_X1 U1550 ( .B1(n19329), .B2(n20304), .C1(n5566), .C2(n20311), .A(
        n2004), .ZN(n2003) );
  OAI221_X1 U1551 ( .B1(n19103), .B2(n1853), .C1(n8482), .C2(n20292), .A(n2005), .ZN(n2002) );
  NOR4_X1 U1552 ( .A1(n1925), .A2(n1926), .A3(n1927), .A4(n1928), .ZN(n1924)
         );
  OAI221_X1 U1553 ( .B1(n8687), .B2(n20234), .C1(n19426), .C2(n20236), .A(
        n1934), .ZN(n1925) );
  OAI221_X1 U1554 ( .B1(n19104), .B2(n1853), .C1(n8483), .C2(n20289), .A(n1930), .ZN(n1927) );
  OAI221_X1 U1555 ( .B1(n19330), .B2(n20300), .C1(n5569), .C2(n20308), .A(
        n1929), .ZN(n1928) );
  NOR4_X1 U1556 ( .A1(n5690), .A2(n5691), .A3(n5692), .A4(n5693), .ZN(n5689)
         );
  OAI221_X1 U1557 ( .B1(n4843), .B2(n20092), .C1(n19363), .C2(n20098), .A(
        n5694), .ZN(n5693) );
  OAI221_X1 U1558 ( .B1(n19075), .B2(n20021), .C1(n18947), .C2(n20025), .A(
        n5708), .ZN(n5690) );
  OAI221_X1 U1559 ( .B1(n19011), .B2(n20047), .C1(n19427), .C2(n20050), .A(
        n5704), .ZN(n5691) );
  NOR4_X1 U1560 ( .A1(n5327), .A2(n5328), .A3(n5329), .A4(n5330), .ZN(n5326)
         );
  OAI221_X1 U1561 ( .B1(n4846), .B2(n20093), .C1(n19364), .C2(n20098), .A(
        n5331), .ZN(n5330) );
  OAI221_X1 U1562 ( .B1(n19076), .B2(n20018), .C1(n18950), .C2(n20027), .A(
        n5631), .ZN(n5327) );
  OAI221_X1 U1563 ( .B1(n19012), .B2(n20047), .C1(n19428), .C2(n20056), .A(
        n5333), .ZN(n5328) );
  NOR4_X1 U1564 ( .A1(n5305), .A2(n5306), .A3(n5307), .A4(n5308), .ZN(n5304)
         );
  OAI221_X1 U1565 ( .B1(n4847), .B2(n20094), .C1(n19365), .C2(n20099), .A(
        n5309), .ZN(n5308) );
  OAI221_X1 U1566 ( .B1(n19077), .B2(n20017), .C1(n18951), .C2(n20026), .A(
        n5313), .ZN(n5305) );
  OAI221_X1 U1567 ( .B1(n19013), .B2(n20048), .C1(n19429), .C2(n20051), .A(
        n5311), .ZN(n5306) );
  NOR4_X1 U1568 ( .A1(n4899), .A2(n4900), .A3(n4901), .A4(n4902), .ZN(n4898)
         );
  OAI221_X1 U1569 ( .B1(n4849), .B2(n20094), .C1(n19366), .C2(n20098), .A(
        n4903), .ZN(n4902) );
  OAI221_X1 U1570 ( .B1(n19078), .B2(n20020), .C1(n18953), .C2(n20027), .A(
        n4907), .ZN(n4899) );
  OAI221_X1 U1571 ( .B1(n19014), .B2(n20047), .C1(n19430), .C2(n20052), .A(
        n4905), .ZN(n4900) );
  NOR4_X1 U1572 ( .A1(n4767), .A2(n4768), .A3(n4769), .A4(n4770), .ZN(n4766)
         );
  OAI221_X1 U1573 ( .B1(n4850), .B2(n20095), .C1(n19367), .C2(n20099), .A(
        n4771), .ZN(n4770) );
  OAI221_X1 U1574 ( .B1(n19079), .B2(n20018), .C1(n18954), .C2(n20028), .A(
        n4775), .ZN(n4767) );
  OAI221_X1 U1575 ( .B1(n19015), .B2(n20048), .C1(n19431), .C2(n20053), .A(
        n4773), .ZN(n4768) );
  NOR4_X1 U1576 ( .A1(n4701), .A2(n4702), .A3(n4703), .A4(n4704), .ZN(n4700)
         );
  OAI221_X1 U1577 ( .B1(n4853), .B2(n20092), .C1(n19368), .C2(n20099), .A(
        n4705), .ZN(n4704) );
  OAI221_X1 U1578 ( .B1(n19080), .B2(n20021), .C1(n18957), .C2(n20030), .A(
        n4709), .ZN(n4701) );
  OAI221_X1 U1579 ( .B1(n19016), .B2(n20048), .C1(n19432), .C2(n20055), .A(
        n4707), .ZN(n4702) );
  NOR4_X1 U1580 ( .A1(n4635), .A2(n4636), .A3(n4637), .A4(n4638), .ZN(n4634)
         );
  OAI221_X1 U1581 ( .B1(n4856), .B2(n20097), .C1(n19369), .C2(n20099), .A(
        n4639), .ZN(n4638) );
  OAI221_X1 U1582 ( .B1(n19081), .B2(n20023), .C1(n18960), .C2(n20028), .A(
        n4643), .ZN(n4635) );
  OAI221_X1 U1583 ( .B1(n19017), .B2(n20048), .C1(n19433), .C2(n20053), .A(
        n4641), .ZN(n4636) );
  NOR4_X1 U1584 ( .A1(n4591), .A2(n4592), .A3(n4593), .A4(n4594), .ZN(n4590)
         );
  OAI221_X1 U1585 ( .B1(n4858), .B2(n20095), .C1(n19370), .C2(n20098), .A(
        n4595), .ZN(n4594) );
  OAI221_X1 U1586 ( .B1(n19082), .B2(n20018), .C1(n18962), .C2(n20028), .A(
        n4599), .ZN(n4591) );
  OAI221_X1 U1587 ( .B1(n19018), .B2(n20047), .C1(n19434), .C2(n20053), .A(
        n4597), .ZN(n4592) );
  NOR4_X1 U1588 ( .A1(n4525), .A2(n4526), .A3(n4527), .A4(n4528), .ZN(n4524)
         );
  OAI221_X1 U1589 ( .B1(n4861), .B2(n20092), .C1(n19371), .C2(n20098), .A(
        n4529), .ZN(n4528) );
  OAI221_X1 U1590 ( .B1(n19019), .B2(n20047), .C1(n19435), .C2(n20055), .A(
        n4531), .ZN(n4526) );
  OAI221_X1 U1591 ( .B1(n19083), .B2(n20021), .C1(n18965), .C2(n20030), .A(
        n4533), .ZN(n4525) );
  NOR4_X1 U1592 ( .A1(n4503), .A2(n4504), .A3(n4505), .A4(n4506), .ZN(n4502)
         );
  OAI221_X1 U1593 ( .B1(n4862), .B2(n20093), .C1(n19372), .C2(n20099), .A(
        n4507), .ZN(n4506) );
  OAI221_X1 U1594 ( .B1(n19020), .B2(n20048), .C1(n19436), .C2(n20050), .A(
        n4509), .ZN(n4504) );
  OAI221_X1 U1595 ( .B1(n19084), .B2(n20019), .C1(n18966), .C2(n20025), .A(
        n4511), .ZN(n4503) );
  NOR4_X1 U1596 ( .A1(n4395), .A2(n4460), .A3(n4461), .A4(n4462), .ZN(n3082)
         );
  OAI221_X1 U1597 ( .B1(n4864), .B2(n20093), .C1(n19373), .C2(n20098), .A(
        n4463), .ZN(n4462) );
  OAI221_X1 U1598 ( .B1(n19021), .B2(n20047), .C1(n19437), .C2(n20054), .A(
        n4465), .ZN(n4460) );
  OAI221_X1 U1599 ( .B1(n19085), .B2(n20022), .C1(n18968), .C2(n20029), .A(
        n4467), .ZN(n4395) );
  NOR4_X1 U1600 ( .A1(n2933), .A2(n2934), .A3(n2935), .A4(n2936), .ZN(n2932)
         );
  OAI221_X1 U1601 ( .B1(n4865), .B2(n20094), .C1(n19374), .C2(n20099), .A(
        n2937), .ZN(n2936) );
  OAI221_X1 U1602 ( .B1(n19086), .B2(n20022), .C1(n18969), .C2(n20031), .A(
        n2941), .ZN(n2933) );
  OAI221_X1 U1603 ( .B1(n19022), .B2(n20048), .C1(n19438), .C2(n20056), .A(
        n2939), .ZN(n2934) );
  NOR4_X1 U1604 ( .A1(n2889), .A2(n2890), .A3(n2891), .A4(n2892), .ZN(n2888)
         );
  OAI221_X1 U1605 ( .B1(n4867), .B2(n20094), .C1(n19375), .C2(n20098), .A(
        n2893), .ZN(n2892) );
  OAI221_X1 U1606 ( .B1(n19087), .B2(n20023), .C1(n18971), .C2(n20027), .A(
        n2897), .ZN(n2889) );
  OAI221_X1 U1607 ( .B1(n19023), .B2(n20047), .C1(n19439), .C2(n20054), .A(
        n2895), .ZN(n2890) );
  NOR4_X1 U1608 ( .A1(n2867), .A2(n2868), .A3(n2869), .A4(n2870), .ZN(n2866)
         );
  OAI221_X1 U1609 ( .B1(n4868), .B2(n20095), .C1(n19376), .C2(n20099), .A(
        n2871), .ZN(n2870) );
  OAI221_X1 U1610 ( .B1(n19088), .B2(n20022), .C1(n18972), .C2(n20027), .A(
        n2875), .ZN(n2867) );
  OAI221_X1 U1611 ( .B1(n19024), .B2(n20048), .C1(n19440), .C2(n20056), .A(
        n2873), .ZN(n2868) );
  NOR4_X1 U1612 ( .A1(n2801), .A2(n2802), .A3(n2803), .A4(n2804), .ZN(n2800)
         );
  OAI221_X1 U1613 ( .B1(n4871), .B2(n20092), .C1(n19377), .C2(n20099), .A(
        n2805), .ZN(n2804) );
  OAI221_X1 U1614 ( .B1(n19089), .B2(n20021), .C1(n18975), .C2(n20025), .A(
        n2809), .ZN(n2801) );
  OAI221_X1 U1615 ( .B1(n19025), .B2(n20048), .C1(n19441), .C2(n20050), .A(
        n2807), .ZN(n2802) );
  NOR4_X1 U1616 ( .A1(n2703), .A2(n2704), .A3(n2705), .A4(n2706), .ZN(n2702)
         );
  OAI221_X1 U1617 ( .B1(n4874), .B2(n20097), .C1(n19378), .C2(n20099), .A(
        n2709), .ZN(n2706) );
  OAI221_X1 U1618 ( .B1(n19090), .B2(n20023), .C1(n18978), .C2(n20028), .A(
        n2725), .ZN(n2703) );
  OAI221_X1 U1619 ( .B1(n19026), .B2(n20048), .C1(n19442), .C2(n20053), .A(
        n2719), .ZN(n2704) );
  NOR4_X1 U1620 ( .A1(n5667), .A2(n5668), .A3(n5669), .A4(n5670), .ZN(n5666)
         );
  OAI221_X1 U1621 ( .B1(n4844), .B2(n20093), .C1(n19379), .C2(n20099), .A(
        n5671), .ZN(n5670) );
  OAI221_X1 U1622 ( .B1(n19091), .B2(n20018), .C1(n18948), .C2(n20026), .A(
        n5675), .ZN(n5667) );
  OAI221_X1 U1623 ( .B1(n19027), .B2(n20048), .C1(n19443), .C2(n20051), .A(
        n5673), .ZN(n5668) );
  NOR4_X1 U1624 ( .A1(n4723), .A2(n4724), .A3(n4725), .A4(n4726), .ZN(n4722)
         );
  OAI221_X1 U1625 ( .B1(n4852), .B2(n20097), .C1(n19380), .C2(n20098), .A(
        n4727), .ZN(n4726) );
  OAI221_X1 U1626 ( .B1(n19092), .B2(n20020), .C1(n18956), .C2(n20031), .A(
        n4731), .ZN(n4723) );
  OAI221_X1 U1627 ( .B1(n19028), .B2(n20047), .C1(n19444), .C2(n20052), .A(
        n4729), .ZN(n4724) );
  NOR4_X1 U1628 ( .A1(n4657), .A2(n4658), .A3(n4659), .A4(n4660), .ZN(n4656)
         );
  OAI221_X1 U1629 ( .B1(n4855), .B2(n20096), .C1(n19381), .C2(n20098), .A(
        n4661), .ZN(n4660) );
  OAI221_X1 U1630 ( .B1(n19093), .B2(n20017), .C1(n18959), .C2(n20026), .A(
        n4665), .ZN(n4657) );
  OAI221_X1 U1631 ( .B1(n19029), .B2(n20047), .C1(n19445), .C2(n20051), .A(
        n4663), .ZN(n4658) );
  NOR4_X1 U1632 ( .A1(n4569), .A2(n4570), .A3(n4571), .A4(n4572), .ZN(n4568)
         );
  OAI221_X1 U1633 ( .B1(n4859), .B2(n20096), .C1(n19382), .C2(n20099), .A(
        n4573), .ZN(n4572) );
  OAI221_X1 U1634 ( .B1(n19094), .B2(n20019), .C1(n18963), .C2(n20029), .A(
        n4577), .ZN(n4569) );
  OAI221_X1 U1635 ( .B1(n19030), .B2(n20048), .C1(n19446), .C2(n20054), .A(
        n4575), .ZN(n4570) );
  NOR4_X1 U1636 ( .A1(n2823), .A2(n2824), .A3(n2825), .A4(n2826), .ZN(n2822)
         );
  OAI221_X1 U1637 ( .B1(n4870), .B2(n20097), .C1(n19383), .C2(n20098), .A(
        n2827), .ZN(n2826) );
  OAI221_X1 U1638 ( .B1(n19095), .B2(n20020), .C1(n18974), .C2(n20031), .A(
        n2831), .ZN(n2823) );
  OAI221_X1 U1639 ( .B1(n19031), .B2(n20047), .C1(n19447), .C2(n20052), .A(
        n2829), .ZN(n2824) );
  NOR4_X1 U1640 ( .A1(n2757), .A2(n2758), .A3(n2759), .A4(n2760), .ZN(n2756)
         );
  OAI221_X1 U1641 ( .B1(n4873), .B2(n20096), .C1(n19384), .C2(n20098), .A(
        n2761), .ZN(n2760) );
  OAI221_X1 U1642 ( .B1(n19096), .B2(n20017), .C1(n18977), .C2(n20026), .A(
        n2765), .ZN(n2757) );
  OAI221_X1 U1643 ( .B1(n19032), .B2(n20047), .C1(n19448), .C2(n20051), .A(
        n2763), .ZN(n2758) );
  NOR4_X1 U1644 ( .A1(n5645), .A2(n5646), .A3(n5647), .A4(n5648), .ZN(n5644)
         );
  OAI221_X1 U1645 ( .B1(n4845), .B2(n20092), .C1(n19385), .C2(n2708), .A(n5649), .ZN(n5648) );
  OAI221_X1 U1646 ( .B1(n19097), .B2(n20022), .C1(n18949), .C2(n20030), .A(
        n5653), .ZN(n5645) );
  OAI221_X1 U1647 ( .B1(n19033), .B2(n2717), .C1(n19449), .C2(n20055), .A(
        n5651), .ZN(n5646) );
  NOR4_X1 U1648 ( .A1(n4745), .A2(n4746), .A3(n4747), .A4(n4748), .ZN(n4744)
         );
  OAI221_X1 U1649 ( .B1(n4851), .B2(n20096), .C1(n19386), .C2(n2708), .A(n4749), .ZN(n4748) );
  OAI221_X1 U1650 ( .B1(n19098), .B2(n20019), .C1(n18955), .C2(n20029), .A(
        n4753), .ZN(n4745) );
  OAI221_X1 U1651 ( .B1(n19034), .B2(n2717), .C1(n19450), .C2(n20054), .A(
        n4751), .ZN(n4746) );
  NOR4_X1 U1652 ( .A1(n4679), .A2(n4680), .A3(n4681), .A4(n4682), .ZN(n4678)
         );
  OAI221_X1 U1653 ( .B1(n4854), .B2(n20093), .C1(n19387), .C2(n2708), .A(n4683), .ZN(n4682) );
  OAI221_X1 U1654 ( .B1(n19099), .B2(n20019), .C1(n18958), .C2(n20030), .A(
        n4687), .ZN(n4679) );
  OAI221_X1 U1655 ( .B1(n19035), .B2(n2717), .C1(n19451), .C2(n20055), .A(
        n4685), .ZN(n4680) );
  NOR4_X1 U1656 ( .A1(n4613), .A2(n4614), .A3(n4615), .A4(n4616), .ZN(n4612)
         );
  OAI221_X1 U1657 ( .B1(n4857), .B2(n20094), .C1(n19388), .C2(n2708), .A(n4617), .ZN(n4616) );
  OAI221_X1 U1658 ( .B1(n19100), .B2(n20019), .C1(n18961), .C2(n20027), .A(
        n4621), .ZN(n4613) );
  OAI221_X1 U1659 ( .B1(n19036), .B2(n2717), .C1(n19452), .C2(n20052), .A(
        n4619), .ZN(n4614) );
  NOR4_X1 U1660 ( .A1(n4547), .A2(n4548), .A3(n4549), .A4(n4550), .ZN(n4546)
         );
  OAI221_X1 U1661 ( .B1(n4860), .B2(n20097), .C1(n19389), .C2(n2708), .A(n4551), .ZN(n4550) );
  OAI221_X1 U1662 ( .B1(n19101), .B2(n20020), .C1(n18964), .C2(n20031), .A(
        n4555), .ZN(n4547) );
  OAI221_X1 U1663 ( .B1(n19037), .B2(n2717), .C1(n19453), .C2(n20052), .A(
        n4553), .ZN(n4548) );
  NOR4_X1 U1664 ( .A1(n4481), .A2(n4482), .A3(n4483), .A4(n4484), .ZN(n4480)
         );
  OAI221_X1 U1665 ( .B1(n4863), .B2(n20092), .C1(n19390), .C2(n2708), .A(n4485), .ZN(n4484) );
  OAI221_X1 U1666 ( .B1(n19038), .B2(n2717), .C1(n19454), .C2(n20054), .A(
        n4487), .ZN(n4482) );
  OAI221_X1 U1667 ( .B1(n19102), .B2(n20017), .C1(n18967), .C2(n20029), .A(
        n4489), .ZN(n4481) );
  NOR4_X1 U1668 ( .A1(n2845), .A2(n2846), .A3(n2847), .A4(n2848), .ZN(n2844)
         );
  OAI221_X1 U1669 ( .B1(n4869), .B2(n20096), .C1(n19391), .C2(n2708), .A(n2849), .ZN(n2848) );
  OAI221_X1 U1670 ( .B1(n19103), .B2(n20023), .C1(n18973), .C2(n20029), .A(
        n2853), .ZN(n2845) );
  OAI221_X1 U1671 ( .B1(n19039), .B2(n2717), .C1(n19455), .C2(n20056), .A(
        n2851), .ZN(n2846) );
  NOR4_X1 U1672 ( .A1(n2779), .A2(n2780), .A3(n2781), .A4(n2782), .ZN(n2778)
         );
  OAI221_X1 U1673 ( .B1(n4872), .B2(n20093), .C1(n19392), .C2(n2708), .A(n2783), .ZN(n2782) );
  OAI221_X1 U1674 ( .B1(n19104), .B2(n20020), .C1(n18976), .C2(n20025), .A(
        n2787), .ZN(n2779) );
  OAI221_X1 U1675 ( .B1(n19040), .B2(n2717), .C1(n19456), .C2(n20050), .A(
        n2785), .ZN(n2780) );
  NOR4_X1 U1676 ( .A1(n4934), .A2(n4935), .A3(n4936), .A4(n4937), .ZN(n4920)
         );
  OAI221_X1 U1677 ( .B1(n4848), .B2(n20095), .C1(n19393), .C2(n2708), .A(n4938), .ZN(n4937) );
  OAI221_X1 U1678 ( .B1(n19105), .B2(n20019), .C1(n18952), .C2(n20029), .A(
        n4942), .ZN(n4934) );
  OAI221_X1 U1679 ( .B1(n19041), .B2(n2717), .C1(n19457), .C2(n20054), .A(
        n4940), .ZN(n4935) );
  NOR4_X1 U1680 ( .A1(n2911), .A2(n2912), .A3(n2913), .A4(n2914), .ZN(n2910)
         );
  OAI221_X1 U1681 ( .B1(n4866), .B2(n20095), .C1(n19394), .C2(n2708), .A(n2915), .ZN(n2914) );
  OAI221_X1 U1682 ( .B1(n19106), .B2(n20018), .C1(n18970), .C2(n20031), .A(
        n2919), .ZN(n2911) );
  OAI221_X1 U1683 ( .B1(n19042), .B2(n2717), .C1(n19458), .C2(n20056), .A(
        n2917), .ZN(n2912) );
  AOI222_X1 U1684 ( .A1(n4739), .A2(n20106), .B1(n3135), .B2(n19780), .C1(
        n2696), .C2(n20585), .ZN(n3136) );
  AOI222_X1 U1685 ( .A1(n4695), .A2(n20104), .B1(n3147), .B2(n19780), .C1(
        n2696), .C2(n20591), .ZN(n3148) );
  AOI222_X1 U1686 ( .A1(n4673), .A2(n20104), .B1(n3153), .B2(n19780), .C1(
        n2696), .C2(n20594), .ZN(n3154) );
  AOI222_X1 U1687 ( .A1(n4629), .A2(n20105), .B1(n3165), .B2(n19780), .C1(
        n2696), .C2(n20600), .ZN(n3166) );
  AOI222_X1 U1688 ( .A1(n4607), .A2(n20105), .B1(n3171), .B2(n19780), .C1(
        n2696), .C2(n20603), .ZN(n3172) );
  AOI222_X1 U1689 ( .A1(n4585), .A2(n20104), .B1(n3177), .B2(n19780), .C1(
        n2696), .C2(n20606), .ZN(n3178) );
  AOI222_X1 U1690 ( .A1(n4541), .A2(n20106), .B1(n3189), .B2(n19780), .C1(
        n2696), .C2(n20612), .ZN(n3190) );
  AOI222_X1 U1691 ( .A1(n4519), .A2(n20105), .B1(n3195), .B2(n19780), .C1(
        n2696), .C2(n20615), .ZN(n3196) );
  AOI222_X1 U1692 ( .A1(n4497), .A2(n20104), .B1(n3201), .B2(n19780), .C1(
        n2696), .C2(n20618), .ZN(n3202) );
  AOI222_X1 U1693 ( .A1(n4475), .A2(n20104), .B1(n3207), .B2(n19779), .C1(
        n2696), .C2(n20621), .ZN(n3208) );
  AOI222_X1 U1694 ( .A1(n2949), .A2(n20106), .B1(n3213), .B2(n19779), .C1(
        n2696), .C2(n20624), .ZN(n3214) );
  AOI222_X1 U1695 ( .A1(n2927), .A2(n20105), .B1(n3219), .B2(n19779), .C1(
        n2696), .C2(n20627), .ZN(n3220) );
  AOI222_X1 U1696 ( .A1(n2883), .A2(n20104), .B1(n3231), .B2(n19779), .C1(
        n2696), .C2(n20633), .ZN(n3232) );
  AOI222_X1 U1697 ( .A1(n2861), .A2(n20106), .B1(n3237), .B2(n19779), .C1(
        n2696), .C2(n20636), .ZN(n3238) );
  AOI222_X1 U1698 ( .A1(n2839), .A2(n20106), .B1(n3243), .B2(n19779), .C1(
        n2696), .C2(n20639), .ZN(n3244) );
  AOI222_X1 U1699 ( .A1(n2795), .A2(n20104), .B1(n3255), .B2(n19779), .C1(
        n2696), .C2(n20645), .ZN(n3256) );
  AOI222_X1 U1700 ( .A1(n2773), .A2(n20104), .B1(n3261), .B2(n19779), .C1(
        n2696), .C2(n20648), .ZN(n3262) );
  AOI222_X1 U1701 ( .A1(n20105), .A2(n2694), .B1(n3273), .B2(n19779), .C1(
        n2696), .C2(n20654), .ZN(n3274) );
  AOI222_X1 U1702 ( .A1(n4717), .A2(n20105), .B1(n3141), .B2(n19780), .C1(
        n2696), .C2(n20588), .ZN(n3142) );
  AOI222_X1 U1703 ( .A1(n4651), .A2(n20106), .B1(n3159), .B2(n19780), .C1(
        n2696), .C2(n20597), .ZN(n3160) );
  AOI222_X1 U1704 ( .A1(n4563), .A2(n20106), .B1(n3183), .B2(n19780), .C1(
        n2696), .C2(n20609), .ZN(n3184) );
  AOI222_X1 U1705 ( .A1(n2905), .A2(n20105), .B1(n3225), .B2(n19779), .C1(
        n2696), .C2(n20630), .ZN(n3226) );
  AOI222_X1 U1706 ( .A1(n2817), .A2(n20105), .B1(n3249), .B2(n19779), .C1(
        n2696), .C2(n20642), .ZN(n3250) );
  AOI222_X1 U1707 ( .A1(n2751), .A2(n20106), .B1(n3267), .B2(n19779), .C1(
        n2696), .C2(n20651), .ZN(n3268) );
  AOI222_X1 U1708 ( .A1(n5683), .A2(n20105), .B1(n3087), .B2(n19781), .C1(
        n2696), .C2(n20561), .ZN(n3088) );
  AOI222_X1 U1709 ( .A1(n5639), .A2(n20104), .B1(n3099), .B2(n19781), .C1(
        n2696), .C2(n20567), .ZN(n3100) );
  AOI222_X1 U1710 ( .A1(n5321), .A2(n20106), .B1(n3105), .B2(n19781), .C1(
        n2696), .C2(n20570), .ZN(n3106) );
  AOI222_X1 U1711 ( .A1(n4950), .A2(n20105), .B1(n3111), .B2(n19781), .C1(
        n2696), .C2(n20573), .ZN(n3112) );
  AOI222_X1 U1712 ( .A1(n4879), .A2(n20104), .B1(n3123), .B2(n19781), .C1(
        n2696), .C2(n20579), .ZN(n3124) );
  AOI222_X1 U1713 ( .A1(n4761), .A2(n20106), .B1(n3129), .B2(n19781), .C1(
        n2696), .C2(n20582), .ZN(n3130) );
  AOI222_X1 U1714 ( .A1(n5661), .A2(n20104), .B1(n3093), .B2(n19781), .C1(
        n2696), .C2(n20564), .ZN(n3094) );
  AOI222_X1 U1715 ( .A1(n4915), .A2(n20105), .B1(n3117), .B2(n19781), .C1(
        n2696), .C2(n20576), .ZN(n3118) );
  AOI222_X1 U1716 ( .A1(n2644), .A2(n20318), .B1(n3277), .B2(n20669), .C1(
        n1837), .C2(n20561), .ZN(n3278) );
  AOI222_X1 U1717 ( .A1(n2619), .A2(n20317), .B1(n3282), .B2(n20669), .C1(
        n1837), .C2(n20564), .ZN(n3283) );
  AOI222_X1 U1718 ( .A1(n2594), .A2(n20317), .B1(n3287), .B2(n20669), .C1(
        n1837), .C2(n20567), .ZN(n3288) );
  AOI222_X1 U1719 ( .A1(n2569), .A2(n20319), .B1(n3292), .B2(n20669), .C1(
        n1837), .C2(n20570), .ZN(n3293) );
  AOI222_X1 U1720 ( .A1(n2544), .A2(n20318), .B1(n3297), .B2(n20669), .C1(
        n1837), .C2(n20573), .ZN(n3298) );
  AOI222_X1 U1721 ( .A1(n2519), .A2(n20318), .B1(n3302), .B2(n20669), .C1(
        n1837), .C2(n20576), .ZN(n3303) );
  AOI222_X1 U1722 ( .A1(n2494), .A2(n20317), .B1(n3307), .B2(n20669), .C1(
        n1837), .C2(n20579), .ZN(n3308) );
  AOI222_X1 U1723 ( .A1(n2469), .A2(n20319), .B1(n3312), .B2(n20669), .C1(
        n1837), .C2(n20582), .ZN(n3313) );
  AOI222_X1 U1724 ( .A1(n2444), .A2(n20319), .B1(n3317), .B2(n20670), .C1(
        n1837), .C2(n20585), .ZN(n3318) );
  AOI222_X1 U1725 ( .A1(n2419), .A2(n20318), .B1(n3322), .B2(n20670), .C1(
        n1837), .C2(n20588), .ZN(n3323) );
  AOI222_X1 U1726 ( .A1(n2394), .A2(n20317), .B1(n3327), .B2(n20670), .C1(
        n1837), .C2(n20591), .ZN(n3328) );
  AOI222_X1 U1727 ( .A1(n2369), .A2(n20317), .B1(n3332), .B2(n20670), .C1(
        n1837), .C2(n20594), .ZN(n3333) );
  AOI222_X1 U1728 ( .A1(n2344), .A2(n20319), .B1(n3337), .B2(n20670), .C1(
        n1837), .C2(n20597), .ZN(n3338) );
  AOI222_X1 U1729 ( .A1(n2319), .A2(n20318), .B1(n3342), .B2(n20670), .C1(
        n1837), .C2(n20600), .ZN(n3343) );
  AOI222_X1 U1730 ( .A1(n2294), .A2(n20318), .B1(n3347), .B2(n20670), .C1(
        n1837), .C2(n20603), .ZN(n3348) );
  AOI222_X1 U1731 ( .A1(n2269), .A2(n20317), .B1(n3352), .B2(n20670), .C1(
        n1837), .C2(n20606), .ZN(n3353) );
  AOI222_X1 U1732 ( .A1(n2244), .A2(n20319), .B1(n3357), .B2(n20670), .C1(
        n1837), .C2(n20609), .ZN(n3358) );
  AOI222_X1 U1733 ( .A1(n2219), .A2(n20319), .B1(n3362), .B2(n20670), .C1(
        n1837), .C2(n20612), .ZN(n3363) );
  AOI222_X1 U1734 ( .A1(n2194), .A2(n20318), .B1(n3367), .B2(n20670), .C1(
        n1837), .C2(n20615), .ZN(n3368) );
  AOI222_X1 U1735 ( .A1(n2169), .A2(n20317), .B1(n3372), .B2(n20670), .C1(
        n1837), .C2(n20618), .ZN(n3373) );
  AOI222_X1 U1736 ( .A1(n2144), .A2(n20317), .B1(n3377), .B2(n20669), .C1(
        n1837), .C2(n20621), .ZN(n3378) );
  AOI222_X1 U1737 ( .A1(n2119), .A2(n20319), .B1(n3382), .B2(n20669), .C1(
        n1837), .C2(n20624), .ZN(n3383) );
  AOI222_X1 U1738 ( .A1(n2094), .A2(n20318), .B1(n3387), .B2(n20669), .C1(
        n1837), .C2(n20627), .ZN(n3388) );
  AOI222_X1 U1739 ( .A1(n2069), .A2(n20318), .B1(n3392), .B2(n20669), .C1(
        n1837), .C2(n20630), .ZN(n3393) );
  AOI222_X1 U1740 ( .A1(n2044), .A2(n20317), .B1(n3397), .B2(n20669), .C1(
        n1837), .C2(n20633), .ZN(n3398) );
  AOI222_X1 U1741 ( .A1(n2019), .A2(n20319), .B1(n3402), .B2(n20669), .C1(
        n1837), .C2(n20636), .ZN(n3403) );
  AOI222_X1 U1742 ( .A1(n1994), .A2(n20319), .B1(n3407), .B2(n20669), .C1(
        n1837), .C2(n20639), .ZN(n3408) );
  AOI222_X1 U1743 ( .A1(n1969), .A2(n20318), .B1(n3412), .B2(n20669), .C1(
        n1837), .C2(n20642), .ZN(n3413) );
  AOI222_X1 U1744 ( .A1(n1944), .A2(n20317), .B1(n3417), .B2(n20669), .C1(
        n1837), .C2(n20645), .ZN(n3418) );
  AOI222_X1 U1745 ( .A1(n1919), .A2(n20317), .B1(n3422), .B2(n20669), .C1(
        n1837), .C2(n20648), .ZN(n3423) );
  AOI222_X1 U1746 ( .A1(n1894), .A2(n20319), .B1(n3427), .B2(n20669), .C1(
        n1837), .C2(n20651), .ZN(n3428) );
  AOI222_X1 U1747 ( .A1(n20318), .A2(n1835), .B1(n3432), .B2(n20669), .C1(
        n1837), .C2(n20654), .ZN(n3433) );
  AND3_X1 U1748 ( .A1(ADD_WR[0]), .A2(n1260), .A3(n1149), .ZN(n1145) );
  AOI21_X1 U1749 ( .B1(n1146), .B2(n5729), .A(n5730), .ZN(n1440) );
  AND2_X1 U1750 ( .A1(n1150), .A2(n1441), .ZN(n5729) );
  INV_X1 U1751 ( .A(WR), .ZN(n5730) );
  OAI221_X1 U1752 ( .B1(n8454), .B2(n20075), .C1(n5126), .C2(n20081), .A(n5702), .ZN(n5692) );
  AOI22_X1 U1753 ( .A1(n20083), .A2(n5835), .B1(n20085), .B2(n5360), .ZN(n5702) );
  OAI221_X1 U1754 ( .B1(n8459), .B2(n20080), .C1(n5128), .C2(n2713), .A(n5650), 
        .ZN(n5647) );
  AOI22_X1 U1755 ( .A1(n20083), .A2(n5837), .B1(n20085), .B2(n5362), .ZN(n5650) );
  OAI221_X1 U1756 ( .B1(n8456), .B2(n20075), .C1(n5129), .C2(n20081), .A(n5332), .ZN(n5329) );
  AOI22_X1 U1757 ( .A1(n2715), .A2(n5838), .B1(n20086), .B2(n5363), .ZN(n5332)
         );
  OAI221_X1 U1758 ( .B1(n8457), .B2(n20078), .C1(n5130), .C2(n20082), .A(n5310), .ZN(n5307) );
  AOI22_X1 U1759 ( .A1(n20083), .A2(n5839), .B1(n20087), .B2(n5364), .ZN(n5310) );
  OAI221_X1 U1760 ( .B1(n8461), .B2(n20076), .C1(n5132), .C2(n20081), .A(n4904), .ZN(n4901) );
  AOI22_X1 U1761 ( .A1(n20083), .A2(n5841), .B1(n20087), .B2(n5366), .ZN(n4904) );
  OAI221_X1 U1762 ( .B1(n8462), .B2(n20076), .C1(n5133), .C2(n20082), .A(n4772), .ZN(n4769) );
  AOI22_X1 U1763 ( .A1(n2715), .A2(n5842), .B1(n20088), .B2(n5367), .ZN(n4772)
         );
  OAI221_X1 U1764 ( .B1(n8467), .B2(n20079), .C1(n5134), .C2(n2713), .A(n4750), 
        .ZN(n4747) );
  AOI22_X1 U1765 ( .A1(n20083), .A2(n5843), .B1(n20089), .B2(n5368), .ZN(n4750) );
  OAI221_X1 U1766 ( .B1(n8464), .B2(n20077), .C1(n5136), .C2(n20082), .A(n4706), .ZN(n4703) );
  AOI22_X1 U1767 ( .A1(n20083), .A2(n5845), .B1(n20085), .B2(n5370), .ZN(n4706) );
  OAI221_X1 U1768 ( .B1(n8468), .B2(n20078), .C1(n5137), .C2(n2713), .A(n4684), 
        .ZN(n4681) );
  AOI22_X1 U1769 ( .A1(n2715), .A2(n5846), .B1(n20086), .B2(n5371), .ZN(n4684)
         );
  OAI221_X1 U1770 ( .B1(n8466), .B2(n20076), .C1(n5139), .C2(n20082), .A(n4640), .ZN(n4637) );
  AOI22_X1 U1771 ( .A1(n2715), .A2(n5848), .B1(n20090), .B2(n5373), .ZN(n4640)
         );
  OAI221_X1 U1772 ( .B1(n8469), .B2(n20076), .C1(n5140), .C2(n2713), .A(n4618), 
        .ZN(n4615) );
  AOI22_X1 U1773 ( .A1(n20083), .A2(n5849), .B1(n20087), .B2(n5374), .ZN(n4618) );
  OAI221_X1 U1774 ( .B1(n8470), .B2(n20076), .C1(n5141), .C2(n20081), .A(n4596), .ZN(n4593) );
  AOI22_X1 U1775 ( .A1(n2715), .A2(n5850), .B1(n20088), .B2(n5375), .ZN(n4596)
         );
  OAI221_X1 U1776 ( .B1(n8473), .B2(n20078), .C1(n5143), .C2(n2713), .A(n4552), 
        .ZN(n4549) );
  AOI22_X1 U1777 ( .A1(n2715), .A2(n5852), .B1(n20090), .B2(n5377), .ZN(n4552)
         );
  OAI221_X1 U1778 ( .B1(n8472), .B2(n20077), .C1(n5144), .C2(n20081), .A(n4530), .ZN(n4527) );
  AOI22_X1 U1779 ( .A1(n20083), .A2(n5853), .B1(n20085), .B2(n5378), .ZN(n4530) );
  OAI221_X1 U1780 ( .B1(n8458), .B2(n20078), .C1(n5145), .C2(n20082), .A(n4508), .ZN(n4505) );
  AOI22_X1 U1781 ( .A1(n2715), .A2(n5854), .B1(n20086), .B2(n5379), .ZN(n4508)
         );
  OAI221_X1 U1782 ( .B1(n8474), .B2(n20077), .C1(n5146), .C2(n2713), .A(n4486), 
        .ZN(n4483) );
  AOI22_X1 U1783 ( .A1(n20083), .A2(n5855), .B1(n20085), .B2(n5440), .ZN(n4486) );
  OAI221_X1 U1784 ( .B1(n8475), .B2(n20078), .C1(n5147), .C2(n20081), .A(n4464), .ZN(n4461) );
  AOI22_X1 U1785 ( .A1(n2715), .A2(n5856), .B1(n20086), .B2(n5441), .ZN(n4464)
         );
  OAI221_X1 U1786 ( .B1(n8476), .B2(n20079), .C1(n5148), .C2(n20082), .A(n2938), .ZN(n2935) );
  AOI22_X1 U1787 ( .A1(n20083), .A2(n5857), .B1(n20087), .B2(n5442), .ZN(n2938) );
  OAI221_X1 U1788 ( .B1(n8478), .B2(n20080), .C1(n5150), .C2(n20081), .A(n2894), .ZN(n2891) );
  AOI22_X1 U1789 ( .A1(n20083), .A2(n5859), .B1(n20087), .B2(n5444), .ZN(n2894) );
  OAI221_X1 U1790 ( .B1(n8479), .B2(n20079), .C1(n4889), .C2(n20082), .A(n2872), .ZN(n2869) );
  AOI22_X1 U1791 ( .A1(n2715), .A2(n5860), .B1(n20088), .B2(n5445), .ZN(n2872)
         );
  OAI221_X1 U1792 ( .B1(n8482), .B2(n20080), .C1(n4890), .C2(n2713), .A(n2850), 
        .ZN(n2847) );
  AOI22_X1 U1793 ( .A1(n20083), .A2(n5861), .B1(n20089), .B2(n5446), .ZN(n2850) );
  OAI221_X1 U1794 ( .B1(n8481), .B2(n20075), .C1(n4892), .C2(n20082), .A(n2806), .ZN(n2803) );
  AOI22_X1 U1795 ( .A1(n20083), .A2(n5863), .B1(n20085), .B2(n5380), .ZN(n2806) );
  OAI221_X1 U1796 ( .B1(n8483), .B2(n20075), .C1(n4893), .C2(n2713), .A(n2784), 
        .ZN(n2781) );
  AOI22_X1 U1797 ( .A1(n2715), .A2(n5864), .B1(n20086), .B2(n5381), .ZN(n2784)
         );
  OAI221_X1 U1798 ( .B1(n8485), .B2(n20075), .C1(n4895), .C2(n20082), .A(n2714), .ZN(n2705) );
  AOI22_X1 U1799 ( .A1(n2715), .A2(n5866), .B1(n20090), .B2(n5383), .ZN(n2714)
         );
  OAI221_X1 U1800 ( .B1(n8455), .B2(n20075), .C1(n5127), .C2(n20082), .A(n5672), .ZN(n5669) );
  AOI22_X1 U1801 ( .A1(n2715), .A2(n5836), .B1(n20086), .B2(n5361), .ZN(n5672)
         );
  OAI221_X1 U1802 ( .B1(n8460), .B2(n20076), .C1(n5131), .C2(n2713), .A(n4939), 
        .ZN(n4936) );
  AOI22_X1 U1803 ( .A1(n2715), .A2(n5840), .B1(n20088), .B2(n5365), .ZN(n4939)
         );
  OAI221_X1 U1804 ( .B1(n8463), .B2(n20077), .C1(n5135), .C2(n20081), .A(n4728), .ZN(n4725) );
  AOI22_X1 U1805 ( .A1(n2715), .A2(n5844), .B1(n20090), .B2(n5369), .ZN(n4728)
         );
  OAI221_X1 U1806 ( .B1(n8465), .B2(n20077), .C1(n5138), .C2(n20081), .A(n4662), .ZN(n4659) );
  AOI22_X1 U1807 ( .A1(n20083), .A2(n5847), .B1(n20089), .B2(n5372), .ZN(n4662) );
  OAI221_X1 U1808 ( .B1(n8471), .B2(n20080), .C1(n5142), .C2(n20082), .A(n4574), .ZN(n4571) );
  AOI22_X1 U1809 ( .A1(n20083), .A2(n5851), .B1(n20089), .B2(n5376), .ZN(n4574) );
  OAI221_X1 U1810 ( .B1(n8477), .B2(n20079), .C1(n5149), .C2(n2713), .A(n2916), 
        .ZN(n2913) );
  AOI22_X1 U1811 ( .A1(n2715), .A2(n5858), .B1(n20088), .B2(n5443), .ZN(n2916)
         );
  OAI221_X1 U1812 ( .B1(n8480), .B2(n20080), .C1(n4891), .C2(n20081), .A(n2828), .ZN(n2825) );
  AOI22_X1 U1813 ( .A1(n2715), .A2(n5862), .B1(n20090), .B2(n5447), .ZN(n2828)
         );
  OAI221_X1 U1814 ( .B1(n8484), .B2(n20079), .C1(n4894), .C2(n20081), .A(n2762), .ZN(n2759) );
  AOI22_X1 U1815 ( .A1(n20083), .A2(n5865), .B1(n20089), .B2(n5382), .ZN(n2762) );
  OAI221_X1 U1816 ( .B1(n19203), .B2(n20266), .C1(n18947), .C2(n20267), .A(
        n2677), .ZN(n2661) );
  AOI22_X1 U1817 ( .A1(n20270), .A2(n5015), .B1(n20279), .B2(n5404), .ZN(n2677) );
  OAI221_X1 U1818 ( .B1(n19204), .B2(n20264), .C1(n18948), .C2(n20268), .A(
        n2633), .ZN(n2626) );
  AOI22_X1 U1819 ( .A1(n20270), .A2(n5016), .B1(n20279), .B2(n5405), .ZN(n2633) );
  OAI221_X1 U1820 ( .B1(n19205), .B2(n20264), .C1(n18949), .C2(n1861), .A(
        n2608), .ZN(n2601) );
  AOI22_X1 U1821 ( .A1(n20274), .A2(n5037), .B1(n20281), .B2(n5406), .ZN(n2608) );
  OAI221_X1 U1822 ( .B1(n19206), .B2(n20263), .C1(n18950), .C2(n20267), .A(
        n2583), .ZN(n2576) );
  AOI22_X1 U1823 ( .A1(n20271), .A2(n5017), .B1(n20280), .B2(n5407), .ZN(n2583) );
  OAI221_X1 U1824 ( .B1(n19207), .B2(n20260), .C1(n18951), .C2(n20268), .A(
        n2558), .ZN(n2551) );
  AOI22_X1 U1825 ( .A1(n20272), .A2(n5018), .B1(n20282), .B2(n5408), .ZN(n2558) );
  OAI221_X1 U1826 ( .B1(n19208), .B2(n20261), .C1(n18952), .C2(n1861), .A(
        n2533), .ZN(n2526) );
  AOI22_X1 U1827 ( .A1(n20272), .A2(n5038), .B1(n20280), .B2(n5409), .ZN(n2533) );
  OAI221_X1 U1828 ( .B1(n19209), .B2(n20260), .C1(n18953), .C2(n20267), .A(
        n2508), .ZN(n2501) );
  AOI22_X1 U1829 ( .A1(n20273), .A2(n5019), .B1(n20281), .B2(n5410), .ZN(n2508) );
  OAI221_X1 U1830 ( .B1(n19210), .B2(n20260), .C1(n18954), .C2(n20268), .A(
        n2483), .ZN(n2476) );
  AOI22_X1 U1831 ( .A1(n20273), .A2(n5020), .B1(n20284), .B2(n5411), .ZN(n2483) );
  OAI221_X1 U1832 ( .B1(n19211), .B2(n20261), .C1(n18955), .C2(n1861), .A(
        n2458), .ZN(n2451) );
  AOI22_X1 U1833 ( .A1(n20272), .A2(n5039), .B1(n20281), .B2(n5412), .ZN(n2458) );
  OAI221_X1 U1834 ( .B1(n19212), .B2(n20262), .C1(n18956), .C2(n20267), .A(
        n2433), .ZN(n2426) );
  AOI22_X1 U1835 ( .A1(n20274), .A2(n5021), .B1(n20282), .B2(n5413), .ZN(n2433) );
  OAI221_X1 U1836 ( .B1(n19213), .B2(n20264), .C1(n18957), .C2(n20268), .A(
        n2408), .ZN(n2401) );
  AOI22_X1 U1837 ( .A1(n20274), .A2(n5022), .B1(n20281), .B2(n5414), .ZN(n2408) );
  OAI221_X1 U1838 ( .B1(n19214), .B2(n20263), .C1(n18958), .C2(n1861), .A(
        n2383), .ZN(n2376) );
  AOI22_X1 U1839 ( .A1(n20275), .A2(n5040), .B1(n20282), .B2(n5415), .ZN(n2383) );
  OAI221_X1 U1840 ( .B1(n19215), .B2(n20260), .C1(n18959), .C2(n20267), .A(
        n2358), .ZN(n2351) );
  AOI22_X1 U1841 ( .A1(n20275), .A2(n5023), .B1(n20283), .B2(n5603), .ZN(n2358) );
  OAI221_X1 U1842 ( .B1(n19216), .B2(n20262), .C1(n18960), .C2(n20268), .A(
        n2333), .ZN(n2326) );
  AOI22_X1 U1843 ( .A1(n20275), .A2(n5024), .B1(n20283), .B2(n5604), .ZN(n2333) );
  OAI221_X1 U1844 ( .B1(n19217), .B2(n20262), .C1(n18961), .C2(n1861), .A(
        n2308), .ZN(n2301) );
  AOI22_X1 U1845 ( .A1(n20274), .A2(n5041), .B1(n20281), .B2(n5605), .ZN(n2308) );
  OAI221_X1 U1846 ( .B1(n19218), .B2(n20260), .C1(n18962), .C2(n20267), .A(
        n2283), .ZN(n2276) );
  AOI22_X1 U1847 ( .A1(n20275), .A2(n5025), .B1(n20282), .B2(n5606), .ZN(n2283) );
  OAI221_X1 U1848 ( .B1(n19219), .B2(n20261), .C1(n18963), .C2(n20268), .A(
        n2258), .ZN(n2251) );
  AOI22_X1 U1849 ( .A1(n20275), .A2(n5026), .B1(n20283), .B2(n5607), .ZN(n2258) );
  OAI221_X1 U1850 ( .B1(n19220), .B2(n20262), .C1(n18964), .C2(n1861), .A(
        n2233), .ZN(n2226) );
  AOI22_X1 U1851 ( .A1(n20275), .A2(n5042), .B1(n20283), .B2(n5608), .ZN(n2233) );
  OAI221_X1 U1852 ( .B1(n19221), .B2(n20265), .C1(n18965), .C2(n20267), .A(
        n2208), .ZN(n2201) );
  AOI22_X1 U1853 ( .A1(n20276), .A2(n5027), .B1(n20284), .B2(n5609), .ZN(n2208) );
  OAI221_X1 U1854 ( .B1(n19222), .B2(n20263), .C1(n18966), .C2(n20268), .A(
        n2183), .ZN(n2176) );
  AOI22_X1 U1855 ( .A1(n20276), .A2(n5028), .B1(n20284), .B2(n5610), .ZN(n2183) );
  OAI221_X1 U1856 ( .B1(n19223), .B2(n20262), .C1(n18967), .C2(n1861), .A(
        n2158), .ZN(n2151) );
  AOI22_X1 U1857 ( .A1(n20276), .A2(n5043), .B1(n20284), .B2(n5629), .ZN(n2158) );
  OAI221_X1 U1858 ( .B1(n19224), .B2(n20264), .C1(n18968), .C2(n20267), .A(
        n2133), .ZN(n2126) );
  AOI22_X1 U1859 ( .A1(n20276), .A2(n5029), .B1(n20284), .B2(n5630), .ZN(n2133) );
  OAI221_X1 U1860 ( .B1(n19225), .B2(n20265), .C1(n18969), .C2(n20268), .A(
        n2108), .ZN(n2101) );
  AOI22_X1 U1861 ( .A1(n20270), .A2(n5030), .B1(n20279), .B2(n5611), .ZN(n2108) );
  OAI221_X1 U1862 ( .B1(n19226), .B2(n20266), .C1(n18970), .C2(n1861), .A(
        n2083), .ZN(n2076) );
  AOI22_X1 U1863 ( .A1(n20274), .A2(n5044), .B1(n20279), .B2(n5612), .ZN(n2083) );
  OAI221_X1 U1864 ( .B1(n19227), .B2(n20266), .C1(n18971), .C2(n20267), .A(
        n2058), .ZN(n2051) );
  AOI22_X1 U1865 ( .A1(n20270), .A2(n5031), .B1(n20279), .B2(n5613), .ZN(n2058) );
  OAI221_X1 U1866 ( .B1(n19228), .B2(n20264), .C1(n18972), .C2(n20268), .A(
        n2033), .ZN(n2026) );
  AOI22_X1 U1867 ( .A1(n20271), .A2(n5032), .B1(n20280), .B2(n5614), .ZN(n2033) );
  OAI221_X1 U1868 ( .B1(n19229), .B2(n20265), .C1(n18973), .C2(n1861), .A(
        n2008), .ZN(n2001) );
  AOI22_X1 U1869 ( .A1(n20271), .A2(n5045), .B1(n20282), .B2(n5615), .ZN(n2008) );
  OAI221_X1 U1870 ( .B1(n19230), .B2(n20261), .C1(n18974), .C2(n20267), .A(
        n1983), .ZN(n1976) );
  AOI22_X1 U1871 ( .A1(n20272), .A2(n5033), .B1(n20280), .B2(n5616), .ZN(n1983) );
  OAI221_X1 U1872 ( .B1(n19231), .B2(n20263), .C1(n18975), .C2(n20268), .A(
        n1958), .ZN(n1951) );
  AOI22_X1 U1873 ( .A1(n20273), .A2(n5034), .B1(n20279), .B2(n5617), .ZN(n1958) );
  OAI221_X1 U1874 ( .B1(n19232), .B2(n20265), .C1(n18976), .C2(n1861), .A(
        n1933), .ZN(n1926) );
  AOI22_X1 U1875 ( .A1(n20271), .A2(n5046), .B1(n20284), .B2(n5618), .ZN(n1933) );
  OAI221_X1 U1876 ( .B1(n19233), .B2(n20265), .C1(n18977), .C2(n20267), .A(
        n1908), .ZN(n1901) );
  AOI22_X1 U1877 ( .A1(n20273), .A2(n5035), .B1(n20283), .B2(n5619), .ZN(n1908) );
  OAI221_X1 U1878 ( .B1(n19234), .B2(n20266), .C1(n18978), .C2(n20268), .A(
        n1862), .ZN(n1845) );
  AOI22_X1 U1879 ( .A1(n20276), .A2(n5036), .B1(n20281), .B2(n5620), .ZN(n1862) );
  NAND4_X1 U1880 ( .A1(n5723), .A2(n1440), .A3(n5724), .A4(n5725), .ZN(n5684)
         );
  NOR3_X1 U1881 ( .A1(n5726), .A2(n5727), .A3(n5728), .ZN(n5725) );
  OAI22_X1 U1882 ( .A1(n4952), .A2(n20124), .B1(n18883), .B2(n20132), .ZN(
        n2692) );
  OAI22_X1 U1883 ( .A1(n4953), .A2(n20125), .B1(n18884), .B2(n20133), .ZN(
        n2642) );
  OAI22_X1 U1884 ( .A1(n4954), .A2(n20124), .B1(n18885), .B2(n20137), .ZN(
        n2617) );
  OAI22_X1 U1885 ( .A1(n4955), .A2(n20130), .B1(n18886), .B2(n20132), .ZN(
        n2592) );
  OAI22_X1 U1886 ( .A1(n4956), .A2(n20126), .B1(n18887), .B2(n20134), .ZN(
        n2567) );
  OAI22_X1 U1887 ( .A1(n4957), .A2(n20127), .B1(n18888), .B2(n20134), .ZN(
        n2542) );
  OAI22_X1 U1888 ( .A1(n4958), .A2(n20127), .B1(n18889), .B2(n20135), .ZN(
        n2517) );
  OAI22_X1 U1889 ( .A1(n4959), .A2(n20127), .B1(n18890), .B2(n20135), .ZN(
        n2492) );
  OAI22_X1 U1890 ( .A1(n4960), .A2(n20128), .B1(n18891), .B2(n20133), .ZN(
        n2467) );
  OAI22_X1 U1891 ( .A1(n4961), .A2(n20126), .B1(n18892), .B2(n20134), .ZN(
        n2442) );
  OAI22_X1 U1892 ( .A1(n4962), .A2(n20129), .B1(n18893), .B2(n20136), .ZN(
        n2417) );
  OAI22_X1 U1893 ( .A1(n4963), .A2(n20130), .B1(n18894), .B2(n20137), .ZN(
        n2392) );
  OAI22_X1 U1894 ( .A1(n4964), .A2(n20126), .B1(n18895), .B2(n20133), .ZN(
        n2367) );
  OAI22_X1 U1895 ( .A1(n4965), .A2(n20127), .B1(n18896), .B2(n20134), .ZN(
        n2342) );
  OAI22_X1 U1896 ( .A1(n4966), .A2(n20127), .B1(n18897), .B2(n20134), .ZN(
        n2317) );
  OAI22_X1 U1897 ( .A1(n4967), .A2(n20128), .B1(n18898), .B2(n20135), .ZN(
        n2292) );
  OAI22_X1 U1898 ( .A1(n4968), .A2(n20128), .B1(n18899), .B2(n20133), .ZN(
        n2267) );
  OAI22_X1 U1899 ( .A1(n4969), .A2(n20125), .B1(n18900), .B2(n20135), .ZN(
        n2242) );
  OAI22_X1 U1900 ( .A1(n4970), .A2(n20129), .B1(n18901), .B2(n20136), .ZN(
        n2217) );
  OAI22_X1 U1901 ( .A1(n4971), .A2(n20128), .B1(n18902), .B2(n20137), .ZN(
        n2192) );
  OAI22_X1 U1902 ( .A1(n4885), .A2(n20124), .B1(n18903), .B2(n20132), .ZN(
        n1967) );
  OAI22_X1 U1903 ( .A1(n4886), .A2(n20125), .B1(n18904), .B2(n20133), .ZN(
        n1942) );
  OAI22_X1 U1904 ( .A1(n4887), .A2(n20124), .B1(n18905), .B2(n20132), .ZN(
        n1917) );
  OAI22_X1 U1905 ( .A1(n4888), .A2(n20129), .B1(n18906), .B2(n20132), .ZN(
        n1890) );
  OAI22_X1 U1906 ( .A1(n8486), .A2(n20212), .B1(n19267), .B2(n20221), .ZN(
        n2683) );
  OAI22_X1 U1907 ( .A1(n8487), .A2(n20212), .B1(n19268), .B2(n20226), .ZN(
        n2638) );
  OAI22_X1 U1908 ( .A1(n8488), .A2(n20212), .B1(n19269), .B2(n20225), .ZN(
        n2613) );
  OAI22_X1 U1909 ( .A1(n8489), .A2(n20212), .B1(n19270), .B2(n20226), .ZN(
        n2588) );
  OAI22_X1 U1910 ( .A1(n8490), .A2(n20213), .B1(n19271), .B2(n20222), .ZN(
        n2563) );
  OAI22_X1 U1911 ( .A1(n8491), .A2(n20214), .B1(n19272), .B2(n20223), .ZN(
        n2538) );
  OAI22_X1 U1912 ( .A1(n8492), .A2(n20214), .B1(n19273), .B2(n20222), .ZN(
        n2513) );
  OAI22_X1 U1913 ( .A1(n8493), .A2(n20213), .B1(n19274), .B2(n20221), .ZN(
        n2488) );
  OAI22_X1 U1914 ( .A1(n8494), .A2(n20218), .B1(n19275), .B2(n20222), .ZN(
        n2463) );
  OAI22_X1 U1915 ( .A1(n8495), .A2(n20216), .B1(n19276), .B2(n20225), .ZN(
        n2438) );
  OAI22_X1 U1916 ( .A1(n8496), .A2(n20215), .B1(n19277), .B2(n20224), .ZN(
        n2413) );
  OAI22_X1 U1917 ( .A1(n8497), .A2(n20216), .B1(n19278), .B2(n20224), .ZN(
        n2388) );
  OAI22_X1 U1918 ( .A1(n8498), .A2(n20213), .B1(n19279), .B2(n20222), .ZN(
        n2363) );
  OAI22_X1 U1919 ( .A1(n8499), .A2(n20214), .B1(n19280), .B2(n20223), .ZN(
        n2338) );
  OAI22_X1 U1920 ( .A1(n8500), .A2(n20213), .B1(n19281), .B2(n20223), .ZN(
        n2313) );
  OAI22_X1 U1921 ( .A1(n8501), .A2(n20214), .B1(n19282), .B2(n20222), .ZN(
        n2288) );
  OAI22_X1 U1922 ( .A1(n8502), .A2(n20213), .B1(n19283), .B2(n20223), .ZN(
        n2263) );
  OAI22_X1 U1923 ( .A1(n8503), .A2(n20217), .B1(n19284), .B2(n20224), .ZN(
        n2238) );
  OAI22_X1 U1924 ( .A1(n8504), .A2(n20215), .B1(n19285), .B2(n20225), .ZN(
        n2213) );
  OAI22_X1 U1925 ( .A1(n8505), .A2(n20216), .B1(n19286), .B2(n20224), .ZN(
        n2188) );
  OAI22_X1 U1926 ( .A1(n8506), .A2(n20216), .B1(n19287), .B2(n20225), .ZN(
        n2163) );
  OAI22_X1 U1927 ( .A1(n8507), .A2(n20217), .B1(n19288), .B2(n20225), .ZN(
        n2138) );
  OAI22_X1 U1928 ( .A1(n8508), .A2(n20217), .B1(n19289), .B2(n20224), .ZN(
        n2113) );
  OAI22_X1 U1929 ( .A1(n8509), .A2(n20218), .B1(n19290), .B2(n20221), .ZN(
        n2088) );
  OAI22_X1 U1930 ( .A1(n8510), .A2(n20218), .B1(n19291), .B2(n20226), .ZN(
        n2063) );
  OAI22_X1 U1931 ( .A1(n8511), .A2(n20218), .B1(n19292), .B2(n20221), .ZN(
        n2038) );
  OAI22_X1 U1932 ( .A1(n8512), .A2(n20215), .B1(n19293), .B2(n20226), .ZN(
        n2013) );
  OAI22_X1 U1933 ( .A1(n8513), .A2(n20217), .B1(n19294), .B2(n20225), .ZN(
        n1988) );
  OAI22_X1 U1934 ( .A1(n8514), .A2(n20212), .B1(n19295), .B2(n20221), .ZN(
        n1963) );
  OAI22_X1 U1935 ( .A1(n8515), .A2(n20212), .B1(n19296), .B2(n20221), .ZN(
        n1938) );
  OAI22_X1 U1936 ( .A1(n8516), .A2(n20215), .B1(n19297), .B2(n20224), .ZN(
        n1913) );
  OAI22_X1 U1937 ( .A1(n8517), .A2(n20218), .B1(n19298), .B2(n20226), .ZN(
        n1874) );
  AND3_X1 U1938 ( .A1(ADD_WR[3]), .A2(n1437), .A3(n1149), .ZN(n1295) );
  OAI22_X1 U1939 ( .A1(n8454), .A2(n19860), .B1(n20561), .B2(n20535), .ZN(
        n4235) );
  OAI22_X1 U1940 ( .A1(n8455), .A2(n19860), .B1(n20564), .B2(n1190), .ZN(n4236) );
  OAI22_X1 U1941 ( .A1(n8456), .A2(n19860), .B1(n20570), .B2(n20535), .ZN(
        n4238) );
  OAI22_X1 U1942 ( .A1(n8457), .A2(n19860), .B1(n20573), .B2(n1190), .ZN(n4239) );
  OAI22_X1 U1943 ( .A1(n8461), .A2(n19860), .B1(n20579), .B2(n20535), .ZN(
        n4241) );
  OAI22_X1 U1944 ( .A1(n8462), .A2(n19860), .B1(n20582), .B2(n1190), .ZN(n4242) );
  OAI22_X1 U1945 ( .A1(n8463), .A2(n19860), .B1(n20588), .B2(n20535), .ZN(
        n4244) );
  OAI22_X1 U1946 ( .A1(n8464), .A2(n19860), .B1(n20591), .B2(n1190), .ZN(n4245) );
  OAI22_X1 U1947 ( .A1(n8465), .A2(n19861), .B1(n20597), .B2(n20535), .ZN(
        n4247) );
  OAI22_X1 U1948 ( .A1(n8466), .A2(n19861), .B1(n20600), .B2(n1190), .ZN(n4248) );
  OAI22_X1 U1949 ( .A1(n8470), .A2(n19861), .B1(n20606), .B2(n20535), .ZN(
        n4250) );
  OAI22_X1 U1950 ( .A1(n8471), .A2(n19861), .B1(n20609), .B2(n1190), .ZN(n4251) );
  OAI22_X1 U1951 ( .A1(n8472), .A2(n19861), .B1(n20615), .B2(n20535), .ZN(
        n4253) );
  OAI22_X1 U1952 ( .A1(n8458), .A2(n19861), .B1(n20618), .B2(n1190), .ZN(n4254) );
  OAI22_X1 U1953 ( .A1(n8475), .A2(n19861), .B1(n20624), .B2(n20535), .ZN(
        n4256) );
  OAI22_X1 U1954 ( .A1(n8476), .A2(n19861), .B1(n20627), .B2(n1190), .ZN(n4257) );
  OAI22_X1 U1955 ( .A1(n8478), .A2(n19862), .B1(n20633), .B2(n20535), .ZN(
        n4259) );
  OAI22_X1 U1956 ( .A1(n8479), .A2(n19862), .B1(n20636), .B2(n1190), .ZN(n4260) );
  OAI22_X1 U1957 ( .A1(n8480), .A2(n19862), .B1(n20642), .B2(n20535), .ZN(
        n4262) );
  OAI22_X1 U1958 ( .A1(n8481), .A2(n19862), .B1(n20645), .B2(n1190), .ZN(n4263) );
  OAI22_X1 U1959 ( .A1(n8484), .A2(n19862), .B1(n20651), .B2(n20535), .ZN(
        n4265) );
  OAI22_X1 U1960 ( .A1(n8485), .A2(n19862), .B1(n20654), .B2(n1190), .ZN(n4266) );
  OAI22_X1 U1961 ( .A1(n8459), .A2(n19860), .B1(n20567), .B2(n20534), .ZN(
        n4237) );
  OAI22_X1 U1962 ( .A1(n8460), .A2(n19860), .B1(n20576), .B2(n20534), .ZN(
        n4240) );
  OAI22_X1 U1963 ( .A1(n8467), .A2(n19860), .B1(n20585), .B2(n20534), .ZN(
        n4243) );
  OAI22_X1 U1964 ( .A1(n8468), .A2(n19860), .B1(n20594), .B2(n20534), .ZN(
        n4246) );
  OAI22_X1 U1965 ( .A1(n8469), .A2(n19861), .B1(n20603), .B2(n20534), .ZN(
        n4249) );
  OAI22_X1 U1966 ( .A1(n8473), .A2(n19861), .B1(n20612), .B2(n20534), .ZN(
        n4252) );
  OAI22_X1 U1967 ( .A1(n8474), .A2(n19861), .B1(n20621), .B2(n20534), .ZN(
        n4255) );
  OAI22_X1 U1968 ( .A1(n8477), .A2(n19861), .B1(n20630), .B2(n20534), .ZN(
        n4258) );
  OAI22_X1 U1969 ( .A1(n8482), .A2(n19862), .B1(n20639), .B2(n20534), .ZN(
        n4261) );
  OAI22_X1 U1970 ( .A1(n8483), .A2(n19862), .B1(n20648), .B2(n20534), .ZN(
        n4264) );
  OAI22_X1 U1971 ( .A1(n20563), .A2(n19890), .B1(n19857), .B2(n19619), .ZN(
        n4203) );
  OAI22_X1 U1972 ( .A1(n20566), .A2(n19891), .B1(n19857), .B2(n19620), .ZN(
        n4204) );
  OAI22_X1 U1973 ( .A1(n20569), .A2(n19891), .B1(n19857), .B2(n19621), .ZN(
        n4205) );
  OAI22_X1 U1974 ( .A1(n20572), .A2(n19892), .B1(n19857), .B2(n19622), .ZN(
        n4206) );
  OAI22_X1 U1975 ( .A1(n20575), .A2(n19890), .B1(n19857), .B2(n19623), .ZN(
        n4207) );
  OAI22_X1 U1976 ( .A1(n20578), .A2(n19892), .B1(n19857), .B2(n19624), .ZN(
        n4208) );
  OAI22_X1 U1977 ( .A1(n20581), .A2(n19891), .B1(n19857), .B2(n19625), .ZN(
        n4209) );
  OAI22_X1 U1978 ( .A1(n20584), .A2(n19892), .B1(n19857), .B2(n19626), .ZN(
        n4210) );
  OAI22_X1 U1979 ( .A1(n20587), .A2(n19890), .B1(n19857), .B2(n19627), .ZN(
        n4211) );
  OAI22_X1 U1980 ( .A1(n20590), .A2(n19890), .B1(n19857), .B2(n19628), .ZN(
        n4212) );
  OAI22_X1 U1981 ( .A1(n20593), .A2(n19891), .B1(n19857), .B2(n19629), .ZN(
        n4213) );
  OAI22_X1 U1982 ( .A1(n20596), .A2(n19891), .B1(n19857), .B2(n19630), .ZN(
        n4214) );
  OAI22_X1 U1983 ( .A1(n20599), .A2(n19892), .B1(n19858), .B2(n19631), .ZN(
        n4215) );
  OAI22_X1 U1984 ( .A1(n20602), .A2(n19890), .B1(n19858), .B2(n19632), .ZN(
        n4216) );
  OAI22_X1 U1985 ( .A1(n20605), .A2(n19892), .B1(n19858), .B2(n19633), .ZN(
        n4217) );
  OAI22_X1 U1986 ( .A1(n20608), .A2(n19891), .B1(n19858), .B2(n19634), .ZN(
        n4218) );
  OAI22_X1 U1987 ( .A1(n20611), .A2(n19892), .B1(n19858), .B2(n19635), .ZN(
        n4219) );
  OAI22_X1 U1988 ( .A1(n20614), .A2(n19890), .B1(n19858), .B2(n19636), .ZN(
        n4220) );
  OAI22_X1 U1989 ( .A1(n20617), .A2(n19890), .B1(n19858), .B2(n19637), .ZN(
        n4221) );
  OAI22_X1 U1990 ( .A1(n20620), .A2(n19891), .B1(n19858), .B2(n19638), .ZN(
        n4222) );
  OAI22_X1 U1991 ( .A1(n20623), .A2(n19891), .B1(n19858), .B2(n19639), .ZN(
        n4223) );
  OAI22_X1 U1992 ( .A1(n20626), .A2(n19892), .B1(n19858), .B2(n19640), .ZN(
        n4224) );
  OAI22_X1 U1993 ( .A1(n20629), .A2(n19890), .B1(n19858), .B2(n19641), .ZN(
        n4225) );
  OAI22_X1 U1994 ( .A1(n20632), .A2(n19892), .B1(n19858), .B2(n19642), .ZN(
        n4226) );
  NAND4_X1 U1995 ( .A1(n2647), .A2(n1440), .A3(n2648), .A4(n2649), .ZN(n2645)
         );
  NOR3_X1 U1996 ( .A1(n2650), .A2(n2651), .A3(n2652), .ZN(n2649) );
  NAND4_X1 U1997 ( .A1(n5686), .A2(n5687), .A3(n5688), .A4(n5689), .ZN(n5685)
         );
  AOI221_X1 U1998 ( .B1(n19900), .B2(n19171), .C1(n19908), .C2(n5768), .A(
        n5721), .ZN(n5686) );
  AOI221_X1 U1999 ( .B1(n19929), .B2(n4997), .C1(n19937), .C2(n5793), .A(n5719), .ZN(n5687) );
  AOI211_X1 U2000 ( .C1(n19961), .C2(n19139), .A(n5711), .B(n5712), .ZN(n5688)
         );
  NAND4_X1 U2001 ( .A1(n5641), .A2(n5642), .A3(n5643), .A4(n5644), .ZN(n5640)
         );
  AOI221_X1 U2002 ( .B1(n19900), .B2(n19173), .C1(n19905), .C2(n5770), .A(
        n5660), .ZN(n5641) );
  AOI221_X1 U2003 ( .B1(n19930), .B2(n4999), .C1(n19937), .C2(n5795), .A(n5659), .ZN(n5642) );
  AOI211_X1 U2004 ( .C1(n19961), .C2(n19141), .A(n5655), .B(n5656), .ZN(n5643)
         );
  NAND4_X1 U2005 ( .A1(n5323), .A2(n5324), .A3(n5325), .A4(n5326), .ZN(n5322)
         );
  AOI221_X1 U2006 ( .B1(n19897), .B2(n19174), .C1(n19906), .C2(n5771), .A(
        n5638), .ZN(n5323) );
  AOI221_X1 U2007 ( .B1(n19931), .B2(n5000), .C1(n19938), .C2(n5796), .A(n5637), .ZN(n5324) );
  AOI211_X1 U2008 ( .C1(n19962), .C2(n19142), .A(n5633), .B(n5634), .ZN(n5325)
         );
  NAND4_X1 U2009 ( .A1(n4976), .A2(n5302), .A3(n5303), .A4(n5304), .ZN(n4951)
         );
  AOI221_X1 U2010 ( .B1(n19898), .B2(n19175), .C1(n19907), .C2(n5772), .A(
        n5320), .ZN(n4976) );
  AOI221_X1 U2011 ( .B1(n19932), .B2(n5270), .C1(n19939), .C2(n5797), .A(n5319), .ZN(n5302) );
  AOI211_X1 U2012 ( .C1(n19963), .C2(n19143), .A(n5315), .B(n5316), .ZN(n5303)
         );
  NAND4_X1 U2013 ( .A1(n4881), .A2(n4896), .A3(n4897), .A4(n4898), .ZN(n4880)
         );
  AOI221_X1 U2014 ( .B1(n19899), .B2(n19177), .C1(n19906), .C2(n5774), .A(
        n4914), .ZN(n4881) );
  AOI221_X1 U2015 ( .B1(n19930), .B2(n5272), .C1(n19940), .C2(n5799), .A(n4913), .ZN(n4896) );
  AOI211_X1 U2016 ( .C1(n19964), .C2(n19145), .A(n4909), .B(n4910), .ZN(n4897)
         );
  NAND4_X1 U2017 ( .A1(n4763), .A2(n4764), .A3(n4765), .A4(n4766), .ZN(n4762)
         );
  AOI221_X1 U2018 ( .B1(n19900), .B2(n19178), .C1(n19908), .C2(n5775), .A(
        n4878), .ZN(n4763) );
  AOI221_X1 U2019 ( .B1(n19932), .B2(n5273), .C1(n19939), .C2(n5800), .A(n4877), .ZN(n4764) );
  AOI211_X1 U2020 ( .C1(n19964), .C2(n19146), .A(n4777), .B(n4778), .ZN(n4765)
         );
  NAND4_X1 U2021 ( .A1(n4741), .A2(n4742), .A3(n4743), .A4(n4744), .ZN(n4740)
         );
  AOI221_X1 U2022 ( .B1(n19902), .B2(n19179), .C1(n19910), .C2(n5776), .A(
        n4760), .ZN(n4741) );
  AOI221_X1 U2023 ( .B1(n19929), .B2(n5274), .C1(n19940), .C2(n5801), .A(n4759), .ZN(n4742) );
  AOI211_X1 U2024 ( .C1(n19963), .C2(n19147), .A(n4755), .B(n4756), .ZN(n4743)
         );
  NAND4_X1 U2025 ( .A1(n4697), .A2(n4698), .A3(n4699), .A4(n4700), .ZN(n4696)
         );
  AOI221_X1 U2026 ( .B1(n19901), .B2(n19181), .C1(n19911), .C2(n5778), .A(
        n4716), .ZN(n4697) );
  AOI221_X1 U2027 ( .B1(n19933), .B2(n5276), .C1(n19941), .C2(n5803), .A(n4715), .ZN(n4698) );
  AOI211_X1 U2028 ( .C1(n19965), .C2(n19149), .A(n4711), .B(n4712), .ZN(n4699)
         );
  NAND4_X1 U2029 ( .A1(n4675), .A2(n4676), .A3(n4677), .A4(n4678), .ZN(n4674)
         );
  AOI221_X1 U2030 ( .B1(n19901), .B2(n19182), .C1(n19909), .C2(n5779), .A(
        n4694), .ZN(n4675) );
  AOI221_X1 U2031 ( .B1(n19933), .B2(n5277), .C1(n19941), .C2(n5804), .A(n4693), .ZN(n4676) );
  AOI211_X1 U2032 ( .C1(n19965), .C2(n19150), .A(n4689), .B(n4690), .ZN(n4677)
         );
  NAND4_X1 U2033 ( .A1(n4631), .A2(n4632), .A3(n4633), .A4(n4634), .ZN(n4630)
         );
  AOI221_X1 U2034 ( .B1(n19902), .B2(n19184), .C1(n19910), .C2(n5781), .A(
        n4650), .ZN(n4631) );
  AOI221_X1 U2035 ( .B1(n19934), .B2(n5279), .C1(n19942), .C2(n5806), .A(n4649), .ZN(n4632) );
  AOI211_X1 U2036 ( .C1(n19967), .C2(n19152), .A(n4645), .B(n4646), .ZN(n4633)
         );
  NAND4_X1 U2037 ( .A1(n4609), .A2(n4610), .A3(n4611), .A4(n4612), .ZN(n4608)
         );
  AOI221_X1 U2038 ( .B1(n19901), .B2(n19185), .C1(n19907), .C2(n5782), .A(
        n4628), .ZN(n4609) );
  AOI221_X1 U2039 ( .B1(n19933), .B2(n5280), .C1(n19941), .C2(n5807), .A(n4627), .ZN(n4610) );
  AOI211_X1 U2040 ( .C1(n19965), .C2(n19153), .A(n4623), .B(n4624), .ZN(n4611)
         );
  NAND4_X1 U2041 ( .A1(n4587), .A2(n4588), .A3(n4589), .A4(n4590), .ZN(n4586)
         );
  AOI221_X1 U2042 ( .B1(n19901), .B2(n19186), .C1(n19909), .C2(n5783), .A(
        n4606), .ZN(n4587) );
  AOI221_X1 U2043 ( .B1(n19932), .B2(n5281), .C1(n19941), .C2(n5808), .A(n4605), .ZN(n4588) );
  AOI211_X1 U2044 ( .C1(n19965), .C2(n19154), .A(n4601), .B(n4602), .ZN(n4589)
         );
  NAND4_X1 U2045 ( .A1(n4543), .A2(n4544), .A3(n4545), .A4(n4546), .ZN(n4542)
         );
  AOI221_X1 U2046 ( .B1(n19902), .B2(n19188), .C1(n19910), .C2(n5785), .A(
        n4562), .ZN(n4543) );
  AOI221_X1 U2047 ( .B1(n19934), .B2(n5283), .C1(n19942), .C2(n5810), .A(n4561), .ZN(n4544) );
  AOI211_X1 U2048 ( .C1(n19966), .C2(n19156), .A(n4557), .B(n4558), .ZN(n4545)
         );
  NAND4_X1 U2049 ( .A1(n4521), .A2(n4522), .A3(n4523), .A4(n4524), .ZN(n4520)
         );
  AOI221_X1 U2050 ( .B1(n19897), .B2(n19189), .C1(n19911), .C2(n5786), .A(
        n4540), .ZN(n4521) );
  AOI221_X1 U2051 ( .B1(n19935), .B2(n5284), .C1(n19943), .C2(n5731), .A(n4539), .ZN(n4522) );
  AOI211_X1 U2052 ( .C1(n19966), .C2(n19157), .A(n4535), .B(n4536), .ZN(n4523)
         );
  NAND4_X1 U2053 ( .A1(n4499), .A2(n4500), .A3(n4501), .A4(n4502), .ZN(n4498)
         );
  AOI221_X1 U2054 ( .B1(n19903), .B2(n19190), .C1(n19911), .C2(n5787), .A(
        n4518), .ZN(n4499) );
  AOI221_X1 U2055 ( .B1(n19935), .B2(n5285), .C1(n19943), .C2(n5732), .A(n4517), .ZN(n4500) );
  AOI211_X1 U2056 ( .C1(n19967), .C2(n19158), .A(n4513), .B(n4514), .ZN(n4501)
         );
  NAND4_X1 U2057 ( .A1(n4477), .A2(n4478), .A3(n4479), .A4(n4480), .ZN(n4476)
         );
  AOI221_X1 U2058 ( .B1(n19903), .B2(n19191), .C1(n19911), .C2(n5883), .A(
        n4496), .ZN(n4477) );
  AOI221_X1 U2059 ( .B1(n19935), .B2(n5621), .C1(n19943), .C2(n5737), .A(n4495), .ZN(n4478) );
  AOI211_X1 U2060 ( .C1(n19966), .C2(n19159), .A(n4491), .B(n4492), .ZN(n4479)
         );
  NAND4_X1 U2061 ( .A1(n2951), .A2(n2952), .A3(n3081), .A4(n3082), .ZN(n2950)
         );
  AOI221_X1 U2062 ( .B1(n19903), .B2(n19192), .C1(n19911), .C2(n5884), .A(
        n4474), .ZN(n2951) );
  AOI221_X1 U2063 ( .B1(n19935), .B2(n5622), .C1(n19943), .C2(n5738), .A(n4473), .ZN(n2952) );
  AOI211_X1 U2064 ( .C1(n19967), .C2(n19160), .A(n4469), .B(n4470), .ZN(n3081)
         );
  NAND4_X1 U2065 ( .A1(n2929), .A2(n2930), .A3(n2931), .A4(n2932), .ZN(n2928)
         );
  AOI221_X1 U2066 ( .B1(n19899), .B2(n19193), .C1(n19905), .C2(n5885), .A(
        n2948), .ZN(n2929) );
  AOI221_X1 U2067 ( .B1(n19929), .B2(n5623), .C1(n19938), .C2(n5739), .A(n2947), .ZN(n2930) );
  AOI211_X1 U2068 ( .C1(n19961), .C2(n19161), .A(n2943), .B(n2944), .ZN(n2931)
         );
  NAND4_X1 U2069 ( .A1(n2885), .A2(n2886), .A3(n2887), .A4(n2888), .ZN(n2884)
         );
  AOI221_X1 U2070 ( .B1(n19897), .B2(n19195), .C1(n19905), .C2(n5886), .A(
        n2904), .ZN(n2885) );
  AOI221_X1 U2071 ( .B1(n19930), .B2(n5625), .C1(n19937), .C2(n5741), .A(n2903), .ZN(n2886) );
  AOI211_X1 U2072 ( .C1(n19966), .C2(n19163), .A(n2899), .B(n2900), .ZN(n2887)
         );
  NAND4_X1 U2073 ( .A1(n2863), .A2(n2864), .A3(n2865), .A4(n2866), .ZN(n2862)
         );
  AOI221_X1 U2074 ( .B1(n19897), .B2(n19196), .C1(n19906), .C2(n5887), .A(
        n2882), .ZN(n2863) );
  AOI221_X1 U2075 ( .B1(n19931), .B2(n5626), .C1(n19938), .C2(n5742), .A(n2881), .ZN(n2864) );
  AOI211_X1 U2076 ( .C1(n19962), .C2(n19164), .A(n2877), .B(n2878), .ZN(n2865)
         );
  NAND4_X1 U2077 ( .A1(n2841), .A2(n2842), .A3(n2843), .A4(n2844), .ZN(n2840)
         );
  AOI221_X1 U2078 ( .B1(n19898), .B2(n19197), .C1(n19907), .C2(n5888), .A(
        n2860), .ZN(n2841) );
  AOI221_X1 U2079 ( .B1(n19932), .B2(n5627), .C1(n19939), .C2(n5743), .A(n2859), .ZN(n2842) );
  AOI211_X1 U2080 ( .C1(n19963), .C2(n19165), .A(n2855), .B(n2856), .ZN(n2843)
         );
  NAND4_X1 U2081 ( .A1(n2797), .A2(n2798), .A3(n2799), .A4(n2800), .ZN(n2796)
         );
  AOI221_X1 U2082 ( .B1(n19899), .B2(n19199), .C1(n19907), .C2(n5788), .A(
        n2816), .ZN(n2797) );
  AOI221_X1 U2083 ( .B1(n19930), .B2(n5286), .C1(n19940), .C2(n5733), .A(n2815), .ZN(n2798) );
  AOI211_X1 U2084 ( .C1(n19964), .C2(n19167), .A(n2811), .B(n2812), .ZN(n2799)
         );
  NAND4_X1 U2085 ( .A1(n2775), .A2(n2776), .A3(n2777), .A4(n2778), .ZN(n2774)
         );
  AOI221_X1 U2086 ( .B1(n19900), .B2(n19200), .C1(n19908), .C2(n5789), .A(
        n2794), .ZN(n2775) );
  AOI221_X1 U2087 ( .B1(n19932), .B2(n5287), .C1(n19938), .C2(n5734), .A(n2793), .ZN(n2776) );
  AOI211_X1 U2088 ( .C1(n19962), .C2(n19168), .A(n2789), .B(n2790), .ZN(n2777)
         );
  NAND4_X1 U2089 ( .A1(n2699), .A2(n2700), .A3(n2701), .A4(n2702), .ZN(n2698)
         );
  AOI221_X1 U2090 ( .B1(n19903), .B2(n19202), .C1(n19909), .C2(n5791), .A(
        n2747), .ZN(n2699) );
  AOI221_X1 U2091 ( .B1(n19929), .B2(n5289), .C1(n19941), .C2(n5736), .A(n2742), .ZN(n2700) );
  AOI211_X1 U2092 ( .C1(n2729), .C2(n19170), .A(n2730), .B(n2731), .ZN(n2701)
         );
  NAND4_X1 U2093 ( .A1(n5663), .A2(n5664), .A3(n5665), .A4(n5666), .ZN(n5662)
         );
  AOI221_X1 U2094 ( .B1(n19900), .B2(n19172), .C1(n19908), .C2(n5769), .A(
        n5682), .ZN(n5663) );
  AOI221_X1 U2095 ( .B1(n19930), .B2(n4998), .C1(n19937), .C2(n5794), .A(n5681), .ZN(n5664) );
  AOI211_X1 U2096 ( .C1(n19961), .C2(n19140), .A(n5677), .B(n5678), .ZN(n5665)
         );
  NAND4_X1 U2097 ( .A1(n4917), .A2(n4918), .A3(n4919), .A4(n4920), .ZN(n4916)
         );
  AOI221_X1 U2098 ( .B1(n19900), .B2(n19176), .C1(n19906), .C2(n5773), .A(
        n4949), .ZN(n4917) );
  AOI221_X1 U2099 ( .B1(n19932), .B2(n5271), .C1(n19938), .C2(n5798), .A(n4948), .ZN(n4918) );
  AOI211_X1 U2100 ( .C1(n19962), .C2(n19144), .A(n4944), .B(n4945), .ZN(n4919)
         );
  NAND4_X1 U2101 ( .A1(n4719), .A2(n4720), .A3(n4721), .A4(n4722), .ZN(n4718)
         );
  AOI221_X1 U2102 ( .B1(n19899), .B2(n19180), .C1(n19909), .C2(n5777), .A(
        n4738), .ZN(n4719) );
  AOI221_X1 U2103 ( .B1(n19933), .B2(n5275), .C1(n19940), .C2(n5802), .A(n4737), .ZN(n4720) );
  AOI211_X1 U2104 ( .C1(n19965), .C2(n19148), .A(n4733), .B(n4734), .ZN(n4721)
         );
  NAND4_X1 U2105 ( .A1(n4653), .A2(n4654), .A3(n4655), .A4(n4656), .ZN(n4652)
         );
  AOI221_X1 U2106 ( .B1(n19902), .B2(n19183), .C1(n19910), .C2(n5780), .A(
        n4672), .ZN(n4653) );
  AOI221_X1 U2107 ( .B1(n19934), .B2(n5278), .C1(n19942), .C2(n5805), .A(n4671), .ZN(n4654) );
  AOI211_X1 U2108 ( .C1(n19967), .C2(n19151), .A(n4667), .B(n4668), .ZN(n4655)
         );
  NAND4_X1 U2109 ( .A1(n4565), .A2(n4566), .A3(n4567), .A4(n4568), .ZN(n4564)
         );
  AOI221_X1 U2110 ( .B1(n19902), .B2(n19187), .C1(n19906), .C2(n5784), .A(
        n4584), .ZN(n4565) );
  AOI221_X1 U2111 ( .B1(n19934), .B2(n5282), .C1(n19942), .C2(n5809), .A(n4583), .ZN(n4566) );
  AOI211_X1 U2112 ( .C1(n19966), .C2(n19155), .A(n4579), .B(n4580), .ZN(n4567)
         );
  NAND4_X1 U2113 ( .A1(n2907), .A2(n2908), .A3(n2909), .A4(n2910), .ZN(n2906)
         );
  AOI221_X1 U2114 ( .B1(n19898), .B2(n19194), .C1(n19905), .C2(n5889), .A(
        n2926), .ZN(n2907) );
  AOI221_X1 U2115 ( .B1(n19929), .B2(n5624), .C1(n19939), .C2(n5740), .A(n2925), .ZN(n2908) );
  AOI211_X1 U2116 ( .C1(n19961), .C2(n19162), .A(n2921), .B(n2922), .ZN(n2909)
         );
  NAND4_X1 U2117 ( .A1(n2819), .A2(n2820), .A3(n2821), .A4(n2822), .ZN(n2818)
         );
  AOI221_X1 U2118 ( .B1(n19901), .B2(n19198), .C1(n19907), .C2(n5890), .A(
        n2838), .ZN(n2819) );
  AOI221_X1 U2119 ( .B1(n19931), .B2(n5628), .C1(n19939), .C2(n5744), .A(n2837), .ZN(n2820) );
  AOI211_X1 U2120 ( .C1(n19963), .C2(n19166), .A(n2833), .B(n2834), .ZN(n2821)
         );
  NAND4_X1 U2121 ( .A1(n2753), .A2(n2754), .A3(n2755), .A4(n2756), .ZN(n2752)
         );
  AOI221_X1 U2122 ( .B1(n19898), .B2(n19201), .C1(n19909), .C2(n5790), .A(
        n2772), .ZN(n2753) );
  AOI221_X1 U2123 ( .B1(n19931), .B2(n5288), .C1(n19937), .C2(n5735), .A(n2771), .ZN(n2754) );
  AOI211_X1 U2124 ( .C1(n19964), .C2(n19169), .A(n2767), .B(n2768), .ZN(n2755)
         );
  NAND4_X1 U2125 ( .A1(n2656), .A2(n2657), .A3(n2658), .A4(n2659), .ZN(n2655)
         );
  AOI221_X1 U2126 ( .B1(n20109), .B2(n19171), .C1(n20120), .C2(n5768), .A(
        n2692), .ZN(n2656) );
  AOI221_X1 U2127 ( .B1(n5176), .B2(n20140), .C1(n20149), .C2(n4779), .A(n2688), .ZN(n2657) );
  AOI211_X1 U2128 ( .C1(n20172), .C2(n19139), .A(n2682), .B(n2683), .ZN(n2658)
         );
  NAND4_X1 U2129 ( .A1(n2621), .A2(n2622), .A3(n2623), .A4(n2624), .ZN(n2620)
         );
  AOI221_X1 U2130 ( .B1(n20110), .B2(n19172), .C1(n20116), .C2(n5769), .A(
        n2642), .ZN(n2621) );
  AOI221_X1 U2131 ( .B1(n5177), .B2(n20141), .C1(n20150), .C2(n4780), .A(n2640), .ZN(n2622) );
  AOI211_X1 U2132 ( .C1(n20172), .C2(n19140), .A(n2637), .B(n2638), .ZN(n2623)
         );
  NAND4_X1 U2133 ( .A1(n2596), .A2(n2597), .A3(n2598), .A4(n2599), .ZN(n2595)
         );
  AOI221_X1 U2134 ( .B1(n20109), .B2(n19173), .C1(n20117), .C2(n5770), .A(
        n2617), .ZN(n2596) );
  AOI221_X1 U2135 ( .B1(n5178), .B2(n20140), .C1(n20150), .C2(n4781), .A(n2615), .ZN(n2597) );
  AOI211_X1 U2136 ( .C1(n20172), .C2(n19141), .A(n2612), .B(n2613), .ZN(n2598)
         );
  NAND4_X1 U2137 ( .A1(n2571), .A2(n2572), .A3(n2573), .A4(n2574), .ZN(n2570)
         );
  AOI221_X1 U2138 ( .B1(n20111), .B2(n19174), .C1(n20116), .C2(n5771), .A(
        n2592), .ZN(n2571) );
  AOI221_X1 U2139 ( .B1(n5179), .B2(n20143), .C1(n20151), .C2(n4782), .A(n2590), .ZN(n2572) );
  AOI211_X1 U2140 ( .C1(n20173), .C2(n19142), .A(n2587), .B(n2588), .ZN(n2573)
         );
  NAND4_X1 U2141 ( .A1(n2546), .A2(n2547), .A3(n2548), .A4(n2549), .ZN(n2545)
         );
  AOI221_X1 U2142 ( .B1(n20111), .B2(n19175), .C1(n20119), .C2(n5772), .A(
        n2567), .ZN(n2546) );
  AOI221_X1 U2143 ( .B1(n5180), .B2(n20142), .C1(n20151), .C2(n4783), .A(n2565), .ZN(n2547) );
  AOI211_X1 U2144 ( .C1(n20173), .C2(n19143), .A(n2562), .B(n2563), .ZN(n2548)
         );
  NAND4_X1 U2145 ( .A1(n2521), .A2(n2522), .A3(n2523), .A4(n2524), .ZN(n2520)
         );
  AOI221_X1 U2146 ( .B1(n20111), .B2(n19176), .C1(n20118), .C2(n5773), .A(
        n2542), .ZN(n2521) );
  AOI221_X1 U2147 ( .B1(n5181), .B2(n20142), .C1(n20151), .C2(n4784), .A(n2540), .ZN(n2522) );
  AOI211_X1 U2148 ( .C1(n20173), .C2(n19144), .A(n2537), .B(n2538), .ZN(n2523)
         );
  NAND4_X1 U2149 ( .A1(n2496), .A2(n2497), .A3(n2498), .A4(n2499), .ZN(n2495)
         );
  AOI221_X1 U2150 ( .B1(n20109), .B2(n19177), .C1(n20118), .C2(n5774), .A(
        n2517), .ZN(n2496) );
  AOI221_X1 U2151 ( .B1(n5182), .B2(n20142), .C1(n20151), .C2(n4785), .A(n2515), .ZN(n2497) );
  AOI211_X1 U2152 ( .C1(n20178), .C2(n19145), .A(n2512), .B(n2513), .ZN(n2498)
         );
  NAND4_X1 U2153 ( .A1(n2471), .A2(n2472), .A3(n2473), .A4(n2474), .ZN(n2470)
         );
  AOI221_X1 U2154 ( .B1(n20113), .B2(n19178), .C1(n20117), .C2(n5775), .A(
        n2492), .ZN(n2471) );
  AOI221_X1 U2155 ( .B1(n5183), .B2(n20144), .C1(n20149), .C2(n4786), .A(n2490), .ZN(n2472) );
  AOI211_X1 U2156 ( .C1(n20174), .C2(n19146), .A(n2487), .B(n2488), .ZN(n2473)
         );
  NAND4_X1 U2157 ( .A1(n2446), .A2(n2447), .A3(n2448), .A4(n2449), .ZN(n2445)
         );
  AOI221_X1 U2158 ( .B1(n20109), .B2(n19179), .C1(n20120), .C2(n5776), .A(
        n2467), .ZN(n2446) );
  AOI221_X1 U2159 ( .B1(n5184), .B2(n20143), .C1(n20150), .C2(n4787), .A(n2465), .ZN(n2447) );
  AOI211_X1 U2160 ( .C1(n20178), .C2(n19147), .A(n2462), .B(n2463), .ZN(n2448)
         );
  NAND4_X1 U2162 ( .A1(n2421), .A2(n2422), .A3(n2423), .A4(n2424), .ZN(n2420)
         );
  AOI221_X1 U2163 ( .B1(n20114), .B2(n19180), .C1(n20119), .C2(n5777), .A(
        n2442), .ZN(n2421) );
  AOI221_X1 U2164 ( .B1(n5185), .B2(n20144), .C1(n20153), .C2(n4788), .A(n2440), .ZN(n2422) );
  AOI211_X1 U2165 ( .C1(n20175), .C2(n19148), .A(n2437), .B(n2438), .ZN(n2423)
         );
  NAND4_X1 U2166 ( .A1(n2396), .A2(n2397), .A3(n2398), .A4(n2399), .ZN(n2395)
         );
  AOI221_X1 U2167 ( .B1(n20112), .B2(n19181), .C1(n20119), .C2(n5778), .A(
        n2417), .ZN(n2396) );
  AOI221_X1 U2168 ( .B1(n5186), .B2(n20145), .C1(n20152), .C2(n4789), .A(n2415), .ZN(n2397) );
  AOI211_X1 U2169 ( .C1(n20175), .C2(n19149), .A(n2412), .B(n2413), .ZN(n2398)
         );
  NAND4_X1 U2170 ( .A1(n2371), .A2(n2372), .A3(n2373), .A4(n2374), .ZN(n2370)
         );
  AOI221_X1 U2171 ( .B1(n20112), .B2(n19182), .C1(n20122), .C2(n5779), .A(
        n2392), .ZN(n2371) );
  AOI221_X1 U2172 ( .B1(n5187), .B2(n20145), .C1(n20152), .C2(n4790), .A(n2390), .ZN(n2372) );
  AOI211_X1 U2173 ( .C1(n20175), .C2(n19150), .A(n2387), .B(n2388), .ZN(n2373)
         );
  NAND4_X1 U2174 ( .A1(n2346), .A2(n2347), .A3(n2348), .A4(n2349), .ZN(n2345)
         );
  AOI221_X1 U2175 ( .B1(n20113), .B2(n19183), .C1(n20120), .C2(n5780), .A(
        n2367), .ZN(n2346) );
  AOI221_X1 U2176 ( .B1(n5188), .B2(n20146), .C1(n20153), .C2(n4791), .A(n2365), .ZN(n2347) );
  AOI211_X1 U2177 ( .C1(n20176), .C2(n19151), .A(n2362), .B(n2363), .ZN(n2348)
         );
  NAND4_X1 U2178 ( .A1(n2321), .A2(n2322), .A3(n2323), .A4(n2324), .ZN(n2320)
         );
  AOI221_X1 U2179 ( .B1(n20114), .B2(n19184), .C1(n20121), .C2(n5781), .A(
        n2342), .ZN(n2321) );
  AOI221_X1 U2180 ( .B1(n5189), .B2(n20142), .C1(n20153), .C2(n4792), .A(n2340), .ZN(n2322) );
  AOI211_X1 U2181 ( .C1(n20177), .C2(n19152), .A(n2337), .B(n2338), .ZN(n2323)
         );
  NAND4_X1 U2182 ( .A1(n2296), .A2(n2297), .A3(n2298), .A4(n2299), .ZN(n2295)
         );
  AOI221_X1 U2183 ( .B1(n20112), .B2(n19185), .C1(n20119), .C2(n5782), .A(
        n2317), .ZN(n2296) );
  AOI221_X1 U2184 ( .B1(n5190), .B2(n20143), .C1(n20152), .C2(n4793), .A(n2315), .ZN(n2297) );
  AOI211_X1 U2185 ( .C1(n20175), .C2(n19153), .A(n2312), .B(n2313), .ZN(n2298)
         );
  NAND4_X1 U2186 ( .A1(n2271), .A2(n2272), .A3(n2273), .A4(n2274), .ZN(n2270)
         );
  AOI221_X1 U2187 ( .B1(n20112), .B2(n19186), .C1(n20120), .C2(n5783), .A(
        n2292), .ZN(n2271) );
  AOI221_X1 U2188 ( .B1(n5191), .B2(n20144), .C1(n20152), .C2(n4794), .A(n2290), .ZN(n2272) );
  AOI211_X1 U2189 ( .C1(n20175), .C2(n19154), .A(n2287), .B(n2288), .ZN(n2273)
         );
  NAND4_X1 U2190 ( .A1(n2246), .A2(n2247), .A3(n2248), .A4(n2249), .ZN(n2245)
         );
  AOI221_X1 U2191 ( .B1(n20113), .B2(n19187), .C1(n20120), .C2(n5784), .A(
        n2267), .ZN(n2246) );
  AOI221_X1 U2192 ( .B1(n5192), .B2(n20145), .C1(n20153), .C2(n4795), .A(n2265), .ZN(n2247) );
  AOI211_X1 U2193 ( .C1(n20176), .C2(n19155), .A(n2262), .B(n2263), .ZN(n2248)
         );
  NAND4_X1 U2194 ( .A1(n2221), .A2(n2222), .A3(n2223), .A4(n2224), .ZN(n2220)
         );
  AOI221_X1 U2195 ( .B1(n20114), .B2(n19188), .C1(n20121), .C2(n5785), .A(
        n2242), .ZN(n2221) );
  AOI221_X1 U2196 ( .B1(n5193), .B2(n20145), .C1(n20153), .C2(n4796), .A(n2240), .ZN(n2222) );
  AOI211_X1 U2197 ( .C1(n20177), .C2(n19156), .A(n2237), .B(n2238), .ZN(n2223)
         );
  NAND4_X1 U2198 ( .A1(n2196), .A2(n2197), .A3(n2198), .A4(n2199), .ZN(n2195)
         );
  AOI221_X1 U2199 ( .B1(n20114), .B2(n19189), .C1(n20122), .C2(n5786), .A(
        n2217), .ZN(n2196) );
  AOI221_X1 U2200 ( .B1(n5194), .B2(n20146), .C1(n20154), .C2(n4797), .A(n2215), .ZN(n2197) );
  AOI211_X1 U2201 ( .C1(n20176), .C2(n19157), .A(n2212), .B(n2213), .ZN(n2198)
         );
  NAND4_X1 U2202 ( .A1(n2171), .A2(n2172), .A3(n2173), .A4(n2174), .ZN(n2170)
         );
  AOI221_X1 U2203 ( .B1(n20113), .B2(n19190), .C1(n20122), .C2(n5787), .A(
        n2192), .ZN(n2171) );
  AOI221_X1 U2204 ( .B1(n5195), .B2(n20146), .C1(n20154), .C2(n4798), .A(n2190), .ZN(n2172) );
  AOI211_X1 U2205 ( .C1(n20177), .C2(n19158), .A(n2187), .B(n2188), .ZN(n2173)
         );
  NAND4_X1 U2206 ( .A1(n2146), .A2(n2147), .A3(n2148), .A4(n2149), .ZN(n2145)
         );
  AOI221_X1 U2207 ( .B1(n20113), .B2(n19191), .C1(n20122), .C2(n5883), .A(
        n2167), .ZN(n2146) );
  AOI221_X1 U2208 ( .B1(n5196), .B2(n20146), .C1(n20154), .C2(n4835), .A(n2165), .ZN(n2147) );
  AOI211_X1 U2209 ( .C1(n20178), .C2(n19159), .A(n2162), .B(n2163), .ZN(n2148)
         );
  NAND4_X1 U2210 ( .A1(n2121), .A2(n2122), .A3(n2123), .A4(n2124), .ZN(n2120)
         );
  AOI221_X1 U2211 ( .B1(n20111), .B2(n19192), .C1(n20122), .C2(n5884), .A(
        n2142), .ZN(n2121) );
  AOI221_X1 U2212 ( .B1(n5197), .B2(n20140), .C1(n20154), .C2(n4836), .A(n2140), .ZN(n2122) );
  AOI211_X1 U2213 ( .C1(n20178), .C2(n19160), .A(n2137), .B(n2138), .ZN(n2123)
         );
  NAND4_X1 U2214 ( .A1(n2096), .A2(n2097), .A3(n2098), .A4(n2099), .ZN(n2095)
         );
  AOI221_X1 U2215 ( .B1(n20109), .B2(n19193), .C1(n20117), .C2(n5885), .A(
        n2117), .ZN(n2096) );
  AOI221_X1 U2216 ( .B1(n5199), .B2(n20144), .C1(n20149), .C2(n4837), .A(n2115), .ZN(n2097) );
  AOI211_X1 U2217 ( .C1(n20172), .C2(n19161), .A(n2112), .B(n2113), .ZN(n2098)
         );
  NAND4_X1 U2218 ( .A1(n2071), .A2(n2072), .A3(n2073), .A4(n2074), .ZN(n2070)
         );
  AOI221_X1 U2219 ( .B1(n20110), .B2(n19194), .C1(n20116), .C2(n5889), .A(
        n2092), .ZN(n2071) );
  AOI221_X1 U2220 ( .B1(n5201), .B2(n20140), .C1(n20150), .C2(n4838), .A(n2090), .ZN(n2072) );
  AOI211_X1 U2221 ( .C1(n20176), .C2(n19162), .A(n2087), .B(n2088), .ZN(n2073)
         );
  NAND4_X1 U2222 ( .A1(n2046), .A2(n2047), .A3(n2048), .A4(n2049), .ZN(n2045)
         );
  AOI221_X1 U2223 ( .B1(n20110), .B2(n19195), .C1(n20117), .C2(n5886), .A(
        n2067), .ZN(n2046) );
  AOI221_X1 U2224 ( .B1(n5203), .B2(n20141), .C1(n20149), .C2(n4839), .A(n2065), .ZN(n2047) );
  AOI211_X1 U2225 ( .C1(n20177), .C2(n19163), .A(n2062), .B(n2063), .ZN(n2048)
         );
  NAND4_X1 U2226 ( .A1(n2021), .A2(n2022), .A3(n2023), .A4(n2024), .ZN(n2020)
         );
  AOI221_X1 U2227 ( .B1(n20114), .B2(n19196), .C1(n20118), .C2(n5887), .A(
        n2042), .ZN(n2021) );
  AOI221_X1 U2228 ( .B1(n5205), .B2(n20140), .C1(n20151), .C2(n4840), .A(n2040), .ZN(n2022) );
  AOI211_X1 U2229 ( .C1(n20173), .C2(n19164), .A(n2037), .B(n2038), .ZN(n2023)
         );
  NAND4_X1 U2230 ( .A1(n1996), .A2(n1997), .A3(n1998), .A4(n1999), .ZN(n1995)
         );
  AOI221_X1 U2231 ( .B1(n20111), .B2(n19197), .C1(n20117), .C2(n5888), .A(
        n2017), .ZN(n1996) );
  AOI221_X1 U2232 ( .B1(n5335), .B2(n20141), .C1(n20149), .C2(n4841), .A(n2015), .ZN(n1997) );
  AOI211_X1 U2233 ( .C1(n20178), .C2(n19165), .A(n2012), .B(n2013), .ZN(n1998)
         );
  NAND4_X1 U2234 ( .A1(n1971), .A2(n1972), .A3(n1973), .A4(n1974), .ZN(n1970)
         );
  AOI221_X1 U2235 ( .B1(n20111), .B2(n19198), .C1(n20118), .C2(n5890), .A(
        n1992), .ZN(n1971) );
  AOI221_X1 U2236 ( .B1(n5337), .B2(n20142), .C1(n20149), .C2(n4842), .A(n1990), .ZN(n1972) );
  AOI211_X1 U2237 ( .C1(n20173), .C2(n19166), .A(n1987), .B(n1988), .ZN(n1973)
         );
  NAND4_X1 U2238 ( .A1(n1946), .A2(n1947), .A3(n1948), .A4(n1949), .ZN(n1945)
         );
  AOI221_X1 U2239 ( .B1(n20112), .B2(n19199), .C1(n20121), .C2(n5788), .A(
        n1967), .ZN(n1946) );
  AOI221_X1 U2240 ( .B1(n5338), .B2(n20141), .C1(n20150), .C2(n4799), .A(n1965), .ZN(n1947) );
  AOI211_X1 U2241 ( .C1(n20174), .C2(n19167), .A(n1962), .B(n1963), .ZN(n1948)
         );
  NAND4_X1 U2242 ( .A1(n1921), .A2(n1922), .A3(n1923), .A4(n1924), .ZN(n1920)
         );
  AOI221_X1 U2243 ( .B1(n20110), .B2(n19200), .C1(n20116), .C2(n5789), .A(
        n1942), .ZN(n1921) );
  AOI221_X1 U2244 ( .B1(n5339), .B2(n20142), .C1(n20151), .C2(n4800), .A(n1940), .ZN(n1922) );
  AOI211_X1 U2245 ( .C1(n20174), .C2(n19168), .A(n1937), .B(n1938), .ZN(n1923)
         );
  NAND4_X1 U2246 ( .A1(n1896), .A2(n1897), .A3(n1898), .A4(n1899), .ZN(n1895)
         );
  AOI221_X1 U2247 ( .B1(n20110), .B2(n19201), .C1(n20121), .C2(n5790), .A(
        n1917), .ZN(n1896) );
  AOI221_X1 U2248 ( .B1(n5340), .B2(n20143), .C1(n20154), .C2(n4801), .A(n1915), .ZN(n1897) );
  AOI211_X1 U2249 ( .C1(n20174), .C2(n19169), .A(n1912), .B(n1913), .ZN(n1898)
         );
  NAND4_X1 U2250 ( .A1(n1840), .A2(n1841), .A3(n1842), .A4(n1843), .ZN(n1839)
         );
  AOI221_X1 U2251 ( .B1(n20112), .B2(n19202), .C1(n20119), .C2(n5791), .A(
        n1890), .ZN(n1840) );
  AOI221_X1 U2252 ( .B1(n1882), .B2(n5341), .C1(n20152), .C2(n4802), .A(n1884), 
        .ZN(n1841) );
  AOI211_X1 U2253 ( .C1(n1871), .C2(n19170), .A(n1873), .B(n1874), .ZN(n1842)
         );
  OAI22_X1 U2254 ( .A1(n20635), .A2(n19891), .B1(n19859), .B2(n19643), .ZN(
        n4227) );
  OAI22_X1 U2255 ( .A1(n20638), .A2(n19892), .B1(n19859), .B2(n19644), .ZN(
        n4228) );
  OAI22_X1 U2256 ( .A1(n20641), .A2(n19890), .B1(n19859), .B2(n19645), .ZN(
        n4229) );
  OAI22_X1 U2257 ( .A1(n20644), .A2(n19890), .B1(n19859), .B2(n19646), .ZN(
        n4230) );
  OAI22_X1 U2258 ( .A1(n20647), .A2(n19891), .B1(n19859), .B2(n19647), .ZN(
        n4231) );
  OAI22_X1 U2259 ( .A1(n20650), .A2(n19891), .B1(n19859), .B2(n19648), .ZN(
        n4232) );
  OAI22_X1 U2260 ( .A1(n20653), .A2(n19892), .B1(n19859), .B2(n19649), .ZN(
        n4233) );
  OAI22_X1 U2261 ( .A1(n20656), .A2(n19890), .B1(n19859), .B2(n19650), .ZN(
        n4234) );
  AOI22_X1 U2262 ( .A1(n20058), .A2(n5290), .B1(n20066), .B2(n19555), .ZN(
        n5704) );
  AOI22_X1 U2263 ( .A1(n20033), .A2(n18979), .B1(n20041), .B2(n19587), .ZN(
        n5708) );
  AOI22_X1 U2264 ( .A1(n20100), .A2(n4921), .B1(n20102), .B2(n4803), .ZN(n5694) );
  AOI22_X1 U2265 ( .A1(n20059), .A2(n5292), .B1(n20067), .B2(n19556), .ZN(
        n5651) );
  AOI22_X1 U2266 ( .A1(n20033), .A2(n18981), .B1(n20041), .B2(n19588), .ZN(
        n5653) );
  AOI22_X1 U2267 ( .A1(n2710), .A2(n4923), .B1(n2711), .B2(n4805), .ZN(n5649)
         );
  AOI22_X1 U2268 ( .A1(n20059), .A2(n5293), .B1(n20068), .B2(n19557), .ZN(
        n5333) );
  AOI22_X1 U2269 ( .A1(n20034), .A2(n18982), .B1(n20042), .B2(n19589), .ZN(
        n5631) );
  AOI22_X1 U2270 ( .A1(n20100), .A2(n4924), .B1(n20102), .B2(n4806), .ZN(n5331) );
  AOI22_X1 U2271 ( .A1(n20058), .A2(n5294), .B1(n20069), .B2(n19558), .ZN(
        n5311) );
  AOI22_X1 U2272 ( .A1(n20034), .A2(n18983), .B1(n20043), .B2(n19590), .ZN(
        n5313) );
  AOI22_X1 U2273 ( .A1(n20101), .A2(n4925), .B1(n20103), .B2(n4807), .ZN(n5309) );
  AOI22_X1 U2274 ( .A1(n20060), .A2(n5296), .B1(n20068), .B2(n19559), .ZN(
        n4905) );
  AOI22_X1 U2275 ( .A1(n20038), .A2(n18985), .B1(n20043), .B2(n19591), .ZN(
        n4907) );
  AOI22_X1 U2276 ( .A1(n20100), .A2(n4927), .B1(n20102), .B2(n4809), .ZN(n4903) );
  AOI22_X1 U2277 ( .A1(n20059), .A2(n5297), .B1(n20067), .B2(n19560), .ZN(
        n4773) );
  AOI22_X1 U2278 ( .A1(n20035), .A2(n18986), .B1(n20044), .B2(n19592), .ZN(
        n4775) );
  AOI22_X1 U2279 ( .A1(n20101), .A2(n4928), .B1(n20103), .B2(n4810), .ZN(n4771) );
  AOI22_X1 U2280 ( .A1(n20063), .A2(n5298), .B1(n20071), .B2(n19561), .ZN(
        n4751) );
  AOI22_X1 U2281 ( .A1(n20034), .A2(n18987), .B1(n20045), .B2(n19593), .ZN(
        n4753) );
  AOI22_X1 U2282 ( .A1(n2710), .A2(n4929), .B1(n2711), .B2(n4811), .ZN(n4749)
         );
  AOI22_X1 U2283 ( .A1(n20061), .A2(n5300), .B1(n20070), .B2(n19562), .ZN(
        n4707) );
  AOI22_X1 U2284 ( .A1(n20036), .A2(n18989), .B1(n20041), .B2(n19594), .ZN(
        n4709) );
  AOI22_X1 U2285 ( .A1(n20101), .A2(n4931), .B1(n20103), .B2(n4813), .ZN(n4705) );
  AOI22_X1 U2286 ( .A1(n20061), .A2(n5301), .B1(n20070), .B2(n19563), .ZN(
        n4685) );
  AOI22_X1 U2287 ( .A1(n20037), .A2(n18990), .B1(n20042), .B2(n19595), .ZN(
        n4687) );
  AOI22_X1 U2288 ( .A1(n2710), .A2(n4932), .B1(n2711), .B2(n4814), .ZN(n4683)
         );
  AOI22_X1 U2289 ( .A1(n20063), .A2(n5385), .B1(n20071), .B2(n19564), .ZN(
        n4641) );
  AOI22_X1 U2290 ( .A1(n20038), .A2(n18992), .B1(n20046), .B2(n19596), .ZN(
        n4643) );
  AOI22_X1 U2291 ( .A1(n20101), .A2(n4978), .B1(n20103), .B2(n4816), .ZN(n4639) );
  AOI22_X1 U2292 ( .A1(n20061), .A2(n5386), .B1(n20070), .B2(n19565), .ZN(
        n4619) );
  AOI22_X1 U2293 ( .A1(n20036), .A2(n18993), .B1(n20043), .B2(n19597), .ZN(
        n4621) );
  AOI22_X1 U2294 ( .A1(n2710), .A2(n4979), .B1(n2711), .B2(n4817), .ZN(n4617)
         );
  AOI22_X1 U2295 ( .A1(n20061), .A2(n5387), .B1(n20070), .B2(n19566), .ZN(
        n4597) );
  AOI22_X1 U2296 ( .A1(n20037), .A2(n18994), .B1(n20044), .B2(n19598), .ZN(
        n4599) );
  AOI22_X1 U2297 ( .A1(n20100), .A2(n4980), .B1(n20102), .B2(n4818), .ZN(n4595) );
  AOI22_X1 U2298 ( .A1(n20063), .A2(n5389), .B1(n20071), .B2(n19567), .ZN(
        n4553) );
  AOI22_X1 U2299 ( .A1(n20038), .A2(n18996), .B1(n20046), .B2(n19599), .ZN(
        n4555) );
  AOI22_X1 U2300 ( .A1(n2710), .A2(n4982), .B1(n2711), .B2(n4820), .ZN(n4551)
         );
  AOI22_X1 U2301 ( .A1(n20037), .A2(n18997), .B1(n20041), .B2(n19600), .ZN(
        n4533) );
  AOI22_X1 U2302 ( .A1(n20063), .A2(n5390), .B1(n20072), .B2(n19568), .ZN(
        n4531) );
  AOI22_X1 U2303 ( .A1(n20100), .A2(n4983), .B1(n20102), .B2(n4821), .ZN(n4529) );
  AOI22_X1 U2304 ( .A1(n20039), .A2(n18998), .B1(n20042), .B2(n19601), .ZN(
        n4511) );
  AOI22_X1 U2305 ( .A1(n20064), .A2(n5391), .B1(n20072), .B2(n19569), .ZN(
        n4509) );
  AOI22_X1 U2306 ( .A1(n20101), .A2(n4984), .B1(n20103), .B2(n4822), .ZN(n4507) );
  AOI22_X1 U2307 ( .A1(n20039), .A2(n18999), .B1(n20041), .B2(n19602), .ZN(
        n4489) );
  AOI22_X1 U2308 ( .A1(n20064), .A2(n5392), .B1(n20072), .B2(n19570), .ZN(
        n4487) );
  AOI22_X1 U2309 ( .A1(n2710), .A2(n4985), .B1(n2711), .B2(n4823), .ZN(n4485)
         );
  AOI22_X1 U2310 ( .A1(n20039), .A2(n19000), .B1(n20042), .B2(n19603), .ZN(
        n4467) );
  AOI22_X1 U2311 ( .A1(n20064), .A2(n5393), .B1(n20072), .B2(n19571), .ZN(
        n4465) );
  AOI22_X1 U2312 ( .A1(n20100), .A2(n4986), .B1(n20102), .B2(n4824), .ZN(n4463) );
  AOI22_X1 U2313 ( .A1(n20058), .A2(n5394), .B1(n20066), .B2(n19572), .ZN(
        n2939) );
  AOI22_X1 U2314 ( .A1(n20033), .A2(n19001), .B1(n20043), .B2(n19604), .ZN(
        n2941) );
  AOI22_X1 U2315 ( .A1(n20101), .A2(n4987), .B1(n20103), .B2(n4825), .ZN(n2937) );
  AOI22_X1 U2316 ( .A1(n20058), .A2(n5396), .B1(n20067), .B2(n19573), .ZN(
        n2895) );
  AOI22_X1 U2317 ( .A1(n20033), .A2(n19003), .B1(n20043), .B2(n19605), .ZN(
        n2897) );
  AOI22_X1 U2318 ( .A1(n20100), .A2(n4989), .B1(n20102), .B2(n4827), .ZN(n2893) );
  AOI22_X1 U2319 ( .A1(n20059), .A2(n5397), .B1(n20068), .B2(n19574), .ZN(
        n2873) );
  AOI22_X1 U2320 ( .A1(n20035), .A2(n19004), .B1(n20044), .B2(n19606), .ZN(
        n2875) );
  AOI22_X1 U2321 ( .A1(n20101), .A2(n4990), .B1(n20103), .B2(n4828), .ZN(n2871) );
  AOI22_X1 U2322 ( .A1(n20058), .A2(n5398), .B1(n20069), .B2(n19575), .ZN(
        n2851) );
  AOI22_X1 U2323 ( .A1(n20034), .A2(n19005), .B1(n20045), .B2(n19607), .ZN(
        n2853) );
  AOI22_X1 U2324 ( .A1(n2710), .A2(n4991), .B1(n2711), .B2(n4829), .ZN(n2849)
         );
  AOI22_X1 U2325 ( .A1(n20060), .A2(n5400), .B1(n20069), .B2(n19576), .ZN(
        n2807) );
  AOI22_X1 U2326 ( .A1(n20039), .A2(n19007), .B1(n20041), .B2(n19608), .ZN(
        n2809) );
  AOI22_X1 U2327 ( .A1(n20101), .A2(n4993), .B1(n20103), .B2(n4831), .ZN(n2805) );
  AOI22_X1 U2328 ( .A1(n20060), .A2(n5401), .B1(n20066), .B2(n19577), .ZN(
        n2785) );
  AOI22_X1 U2329 ( .A1(n20035), .A2(n19008), .B1(n20042), .B2(n19609), .ZN(
        n2787) );
  AOI22_X1 U2330 ( .A1(n2710), .A2(n4994), .B1(n2711), .B2(n4832), .ZN(n2783)
         );
  AOI22_X1 U2331 ( .A1(n20059), .A2(n5403), .B1(n20067), .B2(n19578), .ZN(
        n2719) );
  AOI22_X1 U2332 ( .A1(n20036), .A2(n19010), .B1(n20046), .B2(n19610), .ZN(
        n2725) );
  AOI22_X1 U2333 ( .A1(n20101), .A2(n4996), .B1(n20103), .B2(n4834), .ZN(n2709) );
  AOI22_X1 U2334 ( .A1(n20064), .A2(n5291), .B1(n20068), .B2(n19579), .ZN(
        n5673) );
  AOI22_X1 U2335 ( .A1(n20035), .A2(n18980), .B1(n20042), .B2(n19611), .ZN(
        n5675) );
  AOI22_X1 U2336 ( .A1(n20101), .A2(n4922), .B1(n20103), .B2(n4804), .ZN(n5671) );
  AOI22_X1 U2337 ( .A1(n20062), .A2(n5295), .B1(n20067), .B2(n19580), .ZN(
        n4940) );
  AOI22_X1 U2338 ( .A1(n20038), .A2(n18984), .B1(n20044), .B2(n19612), .ZN(
        n4942) );
  AOI22_X1 U2339 ( .A1(n2710), .A2(n4926), .B1(n2711), .B2(n4808), .ZN(n4938)
         );
  AOI22_X1 U2340 ( .A1(n20060), .A2(n5299), .B1(n20066), .B2(n19581), .ZN(
        n4729) );
  AOI22_X1 U2341 ( .A1(n20035), .A2(n18988), .B1(n20046), .B2(n19613), .ZN(
        n4731) );
  AOI22_X1 U2342 ( .A1(n20100), .A2(n4930), .B1(n20102), .B2(n4812), .ZN(n4727) );
  AOI22_X1 U2343 ( .A1(n20062), .A2(n5384), .B1(n20071), .B2(n19582), .ZN(
        n4663) );
  AOI22_X1 U2344 ( .A1(n20038), .A2(n18991), .B1(n20045), .B2(n19614), .ZN(
        n4665) );
  AOI22_X1 U2345 ( .A1(n20100), .A2(n4933), .B1(n20102), .B2(n4815), .ZN(n4661) );
  AOI22_X1 U2346 ( .A1(n20062), .A2(n5388), .B1(n20069), .B2(n19583), .ZN(
        n4575) );
  AOI22_X1 U2347 ( .A1(n20036), .A2(n18995), .B1(n20045), .B2(n19615), .ZN(
        n4577) );
  AOI22_X1 U2348 ( .A1(n20101), .A2(n4981), .B1(n20103), .B2(n4819), .ZN(n4573) );
  AOI22_X1 U2349 ( .A1(n20064), .A2(n5395), .B1(n20069), .B2(n19584), .ZN(
        n2917) );
  AOI22_X1 U2350 ( .A1(n20037), .A2(n19002), .B1(n20044), .B2(n19616), .ZN(
        n2919) );
  AOI22_X1 U2351 ( .A1(n2710), .A2(n4988), .B1(n2711), .B2(n4826), .ZN(n2915)
         );
  AOI22_X1 U2352 ( .A1(n20062), .A2(n5399), .B1(n20071), .B2(n19585), .ZN(
        n2829) );
  AOI22_X1 U2353 ( .A1(n20037), .A2(n19006), .B1(n20046), .B2(n19617), .ZN(
        n2831) );
  AOI22_X1 U2354 ( .A1(n20100), .A2(n4992), .B1(n20102), .B2(n4830), .ZN(n2827) );
  AOI22_X1 U2355 ( .A1(n20063), .A2(n5402), .B1(n20071), .B2(n19586), .ZN(
        n2763) );
  AOI22_X1 U2356 ( .A1(n20034), .A2(n19009), .B1(n20045), .B2(n19618), .ZN(
        n2765) );
  AOI22_X1 U2357 ( .A1(n20100), .A2(n4995), .B1(n20102), .B2(n4833), .ZN(n2761) );
  AOI22_X1 U2358 ( .A1(n20313), .A2(n4997), .B1(n20315), .B2(n4803), .ZN(n2664) );
  AOI22_X1 U2359 ( .A1(n20294), .A2(n19491), .B1(n20296), .B2(n18979), .ZN(
        n2670) );
  AOI22_X1 U2360 ( .A1(n20248), .A2(n19459), .B1(n20252), .B2(n5047), .ZN(
        n2678) );
  AOI22_X1 U2361 ( .A1(n20314), .A2(n4998), .B1(n20316), .B2(n4804), .ZN(n2629) );
  AOI22_X1 U2362 ( .A1(n20295), .A2(n19492), .B1(n20297), .B2(n18980), .ZN(
        n2630) );
  AOI22_X1 U2363 ( .A1(n20245), .A2(n19460), .B1(n20252), .B2(n5048), .ZN(
        n2634) );
  AOI22_X1 U2364 ( .A1(n1851), .A2(n4999), .B1(n1852), .B2(n4805), .ZN(n2604)
         );
  AOI22_X1 U2365 ( .A1(n1856), .A2(n19493), .B1(n1858), .B2(n18981), .ZN(n2605) );
  AOI22_X1 U2366 ( .A1(n20246), .A2(n19461), .B1(n20252), .B2(n5049), .ZN(
        n2609) );
  AOI22_X1 U2367 ( .A1(n20313), .A2(n5000), .B1(n20315), .B2(n4806), .ZN(n2579) );
  AOI22_X1 U2368 ( .A1(n20294), .A2(n19494), .B1(n20296), .B2(n18982), .ZN(
        n2580) );
  AOI22_X1 U2369 ( .A1(n20244), .A2(n19462), .B1(n20252), .B2(n5050), .ZN(
        n2584) );
  AOI22_X1 U2370 ( .A1(n20314), .A2(n5270), .B1(n20316), .B2(n4807), .ZN(n2554) );
  AOI22_X1 U2371 ( .A1(n20295), .A2(n19495), .B1(n20297), .B2(n18983), .ZN(
        n2555) );
  AOI22_X1 U2372 ( .A1(n20245), .A2(n19463), .B1(n20253), .B2(n5051), .ZN(
        n2559) );
  AOI22_X1 U2373 ( .A1(n1851), .A2(n5271), .B1(n1852), .B2(n4808), .ZN(n2529)
         );
  AOI22_X1 U2374 ( .A1(n1856), .A2(n19496), .B1(n1858), .B2(n18984), .ZN(n2530) );
  AOI22_X1 U2375 ( .A1(n20244), .A2(n19464), .B1(n20253), .B2(n5052), .ZN(
        n2534) );
  AOI22_X1 U2376 ( .A1(n20313), .A2(n5272), .B1(n20315), .B2(n4809), .ZN(n2504) );
  AOI22_X1 U2377 ( .A1(n20294), .A2(n19497), .B1(n20296), .B2(n18985), .ZN(
        n2505) );
  AOI22_X1 U2378 ( .A1(n20246), .A2(n19465), .B1(n20254), .B2(n5053), .ZN(
        n2509) );
  AOI22_X1 U2379 ( .A1(n20314), .A2(n5273), .B1(n20316), .B2(n4810), .ZN(n2479) );
  AOI22_X1 U2380 ( .A1(n20295), .A2(n19498), .B1(n20297), .B2(n18986), .ZN(
        n2480) );
  AOI22_X1 U2381 ( .A1(n20246), .A2(n19466), .B1(n20255), .B2(n5054), .ZN(
        n2484) );
  AOI22_X1 U2382 ( .A1(n1851), .A2(n5274), .B1(n1852), .B2(n4811), .ZN(n2454)
         );
  AOI22_X1 U2383 ( .A1(n1856), .A2(n19499), .B1(n1858), .B2(n18987), .ZN(n2455) );
  AOI22_X1 U2384 ( .A1(n20249), .A2(n19467), .B1(n20254), .B2(n5055), .ZN(
        n2459) );
  AOI22_X1 U2385 ( .A1(n20313), .A2(n5275), .B1(n20315), .B2(n4812), .ZN(n2429) );
  AOI22_X1 U2386 ( .A1(n20294), .A2(n19500), .B1(n20296), .B2(n18988), .ZN(
        n2430) );
  AOI22_X1 U2387 ( .A1(n20246), .A2(n19468), .B1(n20253), .B2(n5056), .ZN(
        n2434) );
  AOI22_X1 U2388 ( .A1(n20314), .A2(n5276), .B1(n20316), .B2(n4813), .ZN(n2404) );
  AOI22_X1 U2389 ( .A1(n20295), .A2(n19501), .B1(n20297), .B2(n18989), .ZN(
        n2405) );
  AOI22_X1 U2390 ( .A1(n20247), .A2(n19469), .B1(n20254), .B2(n5057), .ZN(
        n2409) );
  AOI22_X1 U2391 ( .A1(n1851), .A2(n5277), .B1(n1852), .B2(n4814), .ZN(n2379)
         );
  AOI22_X1 U2392 ( .A1(n1856), .A2(n19502), .B1(n1858), .B2(n18990), .ZN(n2380) );
  AOI22_X1 U2393 ( .A1(n20248), .A2(n19470), .B1(n20256), .B2(n5058), .ZN(
        n2384) );
  AOI22_X1 U2394 ( .A1(n20313), .A2(n5278), .B1(n20315), .B2(n4815), .ZN(n2354) );
  AOI22_X1 U2395 ( .A1(n20294), .A2(n19503), .B1(n20296), .B2(n18991), .ZN(
        n2355) );
  AOI22_X1 U2396 ( .A1(n20249), .A2(n19471), .B1(n20257), .B2(n5059), .ZN(
        n2359) );
  AOI22_X1 U2397 ( .A1(n20314), .A2(n5279), .B1(n20316), .B2(n4816), .ZN(n2329) );
  AOI22_X1 U2398 ( .A1(n20295), .A2(n19504), .B1(n20297), .B2(n18992), .ZN(
        n2330) );
  AOI22_X1 U2399 ( .A1(n20249), .A2(n19472), .B1(n20257), .B2(n5060), .ZN(
        n2334) );
  AOI22_X1 U2400 ( .A1(n1851), .A2(n5280), .B1(n1852), .B2(n4817), .ZN(n2304)
         );
  AOI22_X1 U2401 ( .A1(n1856), .A2(n19505), .B1(n1858), .B2(n18993), .ZN(n2305) );
  AOI22_X1 U2402 ( .A1(n20247), .A2(n19473), .B1(n20255), .B2(n5061), .ZN(
        n2309) );
  AOI22_X1 U2403 ( .A1(n20313), .A2(n5281), .B1(n20315), .B2(n4818), .ZN(n2279) );
  AOI22_X1 U2404 ( .A1(n20294), .A2(n19506), .B1(n20296), .B2(n18994), .ZN(
        n2280) );
  AOI22_X1 U2405 ( .A1(n20248), .A2(n19474), .B1(n20256), .B2(n5062), .ZN(
        n2284) );
  AOI22_X1 U2406 ( .A1(n20314), .A2(n5282), .B1(n20316), .B2(n4819), .ZN(n2254) );
  AOI22_X1 U2407 ( .A1(n20295), .A2(n19507), .B1(n20297), .B2(n18995), .ZN(
        n2255) );
  AOI22_X1 U2408 ( .A1(n20249), .A2(n19475), .B1(n20258), .B2(n5063), .ZN(
        n2259) );
  AOI22_X1 U2409 ( .A1(n1851), .A2(n5283), .B1(n1852), .B2(n4820), .ZN(n2229)
         );
  AOI22_X1 U2410 ( .A1(n1856), .A2(n19508), .B1(n1858), .B2(n18996), .ZN(n2230) );
  AOI22_X1 U2411 ( .A1(n20249), .A2(n19476), .B1(n20257), .B2(n5064), .ZN(
        n2234) );
  AOI22_X1 U2412 ( .A1(n20313), .A2(n5284), .B1(n20315), .B2(n4821), .ZN(n2204) );
  AOI22_X1 U2413 ( .A1(n20294), .A2(n19509), .B1(n20296), .B2(n18997), .ZN(
        n2205) );
  AOI22_X1 U2414 ( .A1(n20250), .A2(n19477), .B1(n20257), .B2(n5065), .ZN(
        n2209) );
  AOI22_X1 U2415 ( .A1(n20314), .A2(n5285), .B1(n20316), .B2(n4822), .ZN(n2179) );
  AOI22_X1 U2416 ( .A1(n20295), .A2(n19510), .B1(n20297), .B2(n18998), .ZN(
        n2180) );
  AOI22_X1 U2417 ( .A1(n20250), .A2(n19478), .B1(n20258), .B2(n5066), .ZN(
        n2184) );
  AOI22_X1 U2418 ( .A1(n1856), .A2(n19511), .B1(n1858), .B2(n18999), .ZN(n2155) );
  AOI22_X1 U2419 ( .A1(n1851), .A2(n5621), .B1(n1852), .B2(n4823), .ZN(n2154)
         );
  AOI22_X1 U2420 ( .A1(n20250), .A2(n19479), .B1(n20258), .B2(n5472), .ZN(
        n2159) );
  AOI22_X1 U2421 ( .A1(n20294), .A2(n19512), .B1(n20296), .B2(n19000), .ZN(
        n2130) );
  AOI22_X1 U2422 ( .A1(n20313), .A2(n5622), .B1(n20315), .B2(n4824), .ZN(n2129) );
  AOI22_X1 U2423 ( .A1(n20250), .A2(n19480), .B1(n20258), .B2(n5473), .ZN(
        n2134) );
  AOI22_X1 U2424 ( .A1(n20295), .A2(n19513), .B1(n20297), .B2(n19001), .ZN(
        n2105) );
  AOI22_X1 U2425 ( .A1(n20314), .A2(n5623), .B1(n20316), .B2(n4825), .ZN(n2104) );
  AOI22_X1 U2426 ( .A1(n20248), .A2(n19481), .B1(n20256), .B2(n5198), .ZN(
        n2109) );
  AOI22_X1 U2427 ( .A1(n1856), .A2(n19514), .B1(n1858), .B2(n19002), .ZN(n2080) );
  AOI22_X1 U2428 ( .A1(n1851), .A2(n5624), .B1(n1852), .B2(n4826), .ZN(n2079)
         );
  AOI22_X1 U2429 ( .A1(n20244), .A2(n19482), .B1(n20252), .B2(n5200), .ZN(
        n2084) );
  AOI22_X1 U2430 ( .A1(n20294), .A2(n19515), .B1(n20296), .B2(n19003), .ZN(
        n2055) );
  AOI22_X1 U2431 ( .A1(n20313), .A2(n5625), .B1(n20315), .B2(n4827), .ZN(n2054) );
  AOI22_X1 U2432 ( .A1(n20248), .A2(n19483), .B1(n20256), .B2(n5202), .ZN(
        n2059) );
  AOI22_X1 U2433 ( .A1(n20295), .A2(n19516), .B1(n20297), .B2(n19004), .ZN(
        n2030) );
  AOI22_X1 U2434 ( .A1(n20314), .A2(n5626), .B1(n20316), .B2(n4828), .ZN(n2029) );
  AOI22_X1 U2435 ( .A1(n20244), .A2(n19484), .B1(n20255), .B2(n5204), .ZN(
        n2034) );
  AOI22_X1 U2436 ( .A1(n1856), .A2(n19517), .B1(n1858), .B2(n19005), .ZN(n2005) );
  AOI22_X1 U2437 ( .A1(n1851), .A2(n5627), .B1(n1852), .B2(n4829), .ZN(n2004)
         );
  AOI22_X1 U2438 ( .A1(n20245), .A2(n19485), .B1(n20253), .B2(n5334), .ZN(
        n2009) );
  AOI22_X1 U2439 ( .A1(n20294), .A2(n19518), .B1(n20296), .B2(n19006), .ZN(
        n1980) );
  AOI22_X1 U2440 ( .A1(n20313), .A2(n5628), .B1(n20315), .B2(n4830), .ZN(n1979) );
  AOI22_X1 U2441 ( .A1(n20245), .A2(n19486), .B1(n20253), .B2(n5336), .ZN(
        n1984) );
  AOI22_X1 U2442 ( .A1(n20314), .A2(n5286), .B1(n20316), .B2(n4831), .ZN(n1954) );
  AOI22_X1 U2443 ( .A1(n20295), .A2(n19519), .B1(n20297), .B2(n19007), .ZN(
        n1955) );
  AOI22_X1 U2444 ( .A1(n20246), .A2(n19487), .B1(n20254), .B2(n5067), .ZN(
        n1959) );
  AOI22_X1 U2445 ( .A1(n1851), .A2(n5287), .B1(n1852), .B2(n4832), .ZN(n1929)
         );
  AOI22_X1 U2446 ( .A1(n1856), .A2(n19520), .B1(n1858), .B2(n19008), .ZN(n1930) );
  AOI22_X1 U2447 ( .A1(n20247), .A2(n19488), .B1(n20255), .B2(n5068), .ZN(
        n1934) );
  AOI22_X1 U2448 ( .A1(n20313), .A2(n5288), .B1(n20315), .B2(n4833), .ZN(n1904) );
  AOI22_X1 U2449 ( .A1(n20294), .A2(n19521), .B1(n20296), .B2(n19009), .ZN(
        n1905) );
  AOI22_X1 U2450 ( .A1(n20250), .A2(n19489), .B1(n20255), .B2(n5069), .ZN(
        n1909) );
  AOI22_X1 U2451 ( .A1(n20314), .A2(n5289), .B1(n20316), .B2(n4834), .ZN(n1850) );
  AOI22_X1 U2452 ( .A1(n20295), .A2(n19522), .B1(n20297), .B2(n19010), .ZN(
        n1855) );
  AOI22_X1 U2453 ( .A1(n20247), .A2(n19490), .B1(n20256), .B2(n5070), .ZN(
        n1867) );
  OAI221_X1 U2454 ( .B1(n19332), .B2(n19969), .C1(n8486), .C2(n19977), .A(
        n5715), .ZN(n5711) );
  AOI22_X1 U2455 ( .A1(n19985), .A2(n5077), .B1(n19993), .B2(n19523), .ZN(
        n5715) );
  OAI221_X1 U2456 ( .B1(n19333), .B2(n19970), .C1(n8488), .C2(n19979), .A(
        n5657), .ZN(n5655) );
  AOI22_X1 U2457 ( .A1(n19986), .A2(n5079), .B1(n19994), .B2(n19524), .ZN(
        n5657) );
  OAI221_X1 U2458 ( .B1(n19334), .B2(n19971), .C1(n8489), .C2(n19980), .A(
        n5635), .ZN(n5633) );
  AOI22_X1 U2459 ( .A1(n19986), .A2(n5080), .B1(n19995), .B2(n19525), .ZN(
        n5635) );
  OAI221_X1 U2460 ( .B1(n19335), .B2(n19970), .C1(n8490), .C2(n19979), .A(
        n5317), .ZN(n5315) );
  AOI22_X1 U2461 ( .A1(n19987), .A2(n5081), .B1(n19996), .B2(n19526), .ZN(
        n5317) );
  OAI221_X1 U2462 ( .B1(n19336), .B2(n19971), .C1(n8492), .C2(n19980), .A(
        n4911), .ZN(n4909) );
  AOI22_X1 U2463 ( .A1(n19988), .A2(n5083), .B1(n19996), .B2(n19527), .ZN(
        n4911) );
  OAI221_X1 U2464 ( .B1(n19337), .B2(n19972), .C1(n8493), .C2(n19981), .A(
        n4875), .ZN(n4777) );
  AOI22_X1 U2465 ( .A1(n19985), .A2(n5084), .B1(n19994), .B2(n19528), .ZN(
        n4875) );
  OAI221_X1 U2466 ( .B1(n19338), .B2(n19970), .C1(n8494), .C2(n19982), .A(
        n4757), .ZN(n4755) );
  AOI22_X1 U2467 ( .A1(n19985), .A2(n5085), .B1(n19998), .B2(n19529), .ZN(
        n4757) );
  OAI221_X1 U2468 ( .B1(n19339), .B2(n19970), .C1(n8496), .C2(n19982), .A(
        n4713), .ZN(n4711) );
  AOI22_X1 U2469 ( .A1(n19989), .A2(n5087), .B1(n19997), .B2(n19530), .ZN(
        n4713) );
  OAI221_X1 U2470 ( .B1(n19340), .B2(n19973), .C1(n8497), .C2(n19982), .A(
        n4691), .ZN(n4689) );
  AOI22_X1 U2471 ( .A1(n19989), .A2(n5088), .B1(n19997), .B2(n19531), .ZN(
        n4691) );
  OAI221_X1 U2472 ( .B1(n19341), .B2(n19972), .C1(n8499), .C2(n19981), .A(
        n4647), .ZN(n4645) );
  AOI22_X1 U2473 ( .A1(n19990), .A2(n5090), .B1(n19998), .B2(n19532), .ZN(
        n4647) );
  OAI221_X1 U2474 ( .B1(n19342), .B2(n19971), .C1(n8500), .C2(n19980), .A(
        n4625), .ZN(n4623) );
  AOI22_X1 U2475 ( .A1(n19989), .A2(n5091), .B1(n19997), .B2(n19533), .ZN(
        n4625) );
  OAI221_X1 U2476 ( .B1(n19343), .B2(n19972), .C1(n8501), .C2(n19981), .A(
        n4603), .ZN(n4601) );
  AOI22_X1 U2477 ( .A1(n19988), .A2(n5092), .B1(n19997), .B2(n19534), .ZN(
        n4603) );
  OAI221_X1 U2478 ( .B1(n19344), .B2(n19970), .C1(n8503), .C2(n19982), .A(
        n4559), .ZN(n4557) );
  AOI22_X1 U2479 ( .A1(n19990), .A2(n5151), .B1(n19998), .B2(n19535), .ZN(
        n4559) );
  OAI221_X1 U2480 ( .B1(n19345), .B2(n19973), .C1(n8504), .C2(n19979), .A(
        n4537), .ZN(n4535) );
  AOI22_X1 U2481 ( .A1(n19991), .A2(n5001), .B1(n19999), .B2(n19536), .ZN(
        n4537) );
  OAI221_X1 U2482 ( .B1(n19346), .B2(n19973), .C1(n8505), .C2(n19982), .A(
        n4515), .ZN(n4513) );
  AOI22_X1 U2483 ( .A1(n19991), .A2(n5002), .B1(n19999), .B2(n19537), .ZN(
        n4515) );
  OAI221_X1 U2484 ( .B1(n19347), .B2(n19974), .C1(n8506), .C2(n19978), .A(
        n4493), .ZN(n4491) );
  AOI22_X1 U2485 ( .A1(n19991), .A2(n5007), .B1(n19999), .B2(n19538), .ZN(
        n4493) );
  OAI221_X1 U2486 ( .B1(n19348), .B2(n19975), .C1(n8507), .C2(n19977), .A(
        n4471), .ZN(n4469) );
  AOI22_X1 U2487 ( .A1(n19991), .A2(n5008), .B1(n19999), .B2(n19539), .ZN(
        n4471) );
  OAI221_X1 U2488 ( .B1(n19349), .B2(n19969), .C1(n8508), .C2(n19983), .A(
        n2945), .ZN(n2943) );
  AOI22_X1 U2489 ( .A1(n19985), .A2(n5009), .B1(n19993), .B2(n19540), .ZN(
        n2945) );
  OAI221_X1 U2490 ( .B1(n19350), .B2(n19974), .C1(n8510), .C2(n19977), .A(
        n2901), .ZN(n2899) );
  AOI22_X1 U2491 ( .A1(n19986), .A2(n5011), .B1(n19994), .B2(n19541), .ZN(
        n2901) );
  OAI221_X1 U2492 ( .B1(n19351), .B2(n19974), .C1(n8511), .C2(n19983), .A(
        n2879), .ZN(n2877) );
  AOI22_X1 U2493 ( .A1(n19990), .A2(n5012), .B1(n19995), .B2(n19542), .ZN(
        n2879) );
  OAI221_X1 U2494 ( .B1(n19352), .B2(n19975), .C1(n8512), .C2(n19983), .A(
        n2857), .ZN(n2855) );
  AOI22_X1 U2495 ( .A1(n19987), .A2(n5013), .B1(n19996), .B2(n19543), .ZN(
        n2857) );
  OAI221_X1 U2496 ( .B1(n19353), .B2(n19969), .C1(n8514), .C2(n19977), .A(
        n2813), .ZN(n2811) );
  AOI22_X1 U2497 ( .A1(n19988), .A2(n5003), .B1(n19995), .B2(n19544), .ZN(
        n2813) );
  OAI221_X1 U2498 ( .B1(n19354), .B2(n19975), .C1(n8515), .C2(n19978), .A(
        n2791), .ZN(n2789) );
  AOI22_X1 U2499 ( .A1(n19986), .A2(n5004), .B1(n19993), .B2(n19545), .ZN(
        n2791) );
  OAI221_X1 U2500 ( .B1(n19331), .B2(n19972), .C1(n8517), .C2(n19981), .A(
        n2736), .ZN(n2730) );
  AOI22_X1 U2501 ( .A1(n19987), .A2(n5006), .B1(n19994), .B2(n19546), .ZN(
        n2736) );
  OAI221_X1 U2502 ( .B1(n19355), .B2(n19969), .C1(n8487), .C2(n19978), .A(
        n5679), .ZN(n5677) );
  AOI22_X1 U2503 ( .A1(n19985), .A2(n5078), .B1(n19996), .B2(n19547), .ZN(
        n5679) );
  OAI221_X1 U2504 ( .B1(n19356), .B2(n19971), .C1(n8491), .C2(n19980), .A(
        n4946), .ZN(n4944) );
  AOI22_X1 U2505 ( .A1(n19988), .A2(n5082), .B1(n19998), .B2(n19548), .ZN(
        n4946) );
  OAI221_X1 U2506 ( .B1(n19357), .B2(n19973), .C1(n8495), .C2(n19979), .A(
        n4735), .ZN(n4733) );
  AOI22_X1 U2507 ( .A1(n19989), .A2(n5086), .B1(n19993), .B2(n19549), .ZN(
        n4735) );
  OAI221_X1 U2508 ( .B1(n19358), .B2(n19970), .C1(n8498), .C2(n19979), .A(
        n4669), .ZN(n4667) );
  AOI22_X1 U2509 ( .A1(n19988), .A2(n5089), .B1(n19995), .B2(n19550), .ZN(
        n4669) );
  OAI221_X1 U2510 ( .B1(n19359), .B2(n19973), .C1(n8502), .C2(n19979), .A(
        n4581), .ZN(n4579) );
  AOI22_X1 U2511 ( .A1(n19990), .A2(n5093), .B1(n19998), .B2(n19551), .ZN(
        n4581) );
  OAI221_X1 U2512 ( .B1(n19360), .B2(n19974), .C1(n8509), .C2(n19983), .A(
        n2923), .ZN(n2921) );
  AOI22_X1 U2513 ( .A1(n19986), .A2(n5010), .B1(n19995), .B2(n19552), .ZN(
        n2923) );
  OAI221_X1 U2514 ( .B1(n19361), .B2(n19975), .C1(n8513), .C2(n19978), .A(
        n2835), .ZN(n2833) );
  AOI22_X1 U2515 ( .A1(n19987), .A2(n5014), .B1(n19998), .B2(n19553), .ZN(
        n2835) );
  OAI221_X1 U2516 ( .B1(n19362), .B2(n19973), .C1(n8516), .C2(n19982), .A(
        n2769), .ZN(n2767) );
  AOI22_X1 U2517 ( .A1(n19990), .A2(n5005), .B1(n19993), .B2(n19554), .ZN(
        n2769) );
  OAI221_X1 U2518 ( .B1(n18915), .B2(n20180), .C1(n19107), .C2(n20193), .A(
        n2686), .ZN(n2682) );
  AOI22_X1 U2519 ( .A1(n20196), .A2(n5360), .B1(n20205), .B2(n5077), .ZN(n2686) );
  OAI221_X1 U2520 ( .B1(n18916), .B2(n20186), .C1(n19108), .C2(n20192), .A(
        n2639), .ZN(n2637) );
  AOI22_X1 U2521 ( .A1(n20202), .A2(n5361), .B1(n20209), .B2(n5078), .ZN(n2639) );
  OAI221_X1 U2522 ( .B1(n18917), .B2(n20186), .C1(n19109), .C2(n20192), .A(
        n2614), .ZN(n2612) );
  AOI22_X1 U2523 ( .A1(n20201), .A2(n5362), .B1(n20210), .B2(n5079), .ZN(n2614) );
  OAI221_X1 U2524 ( .B1(n18918), .B2(n20184), .C1(n19110), .C2(n20193), .A(
        n2589), .ZN(n2587) );
  AOI22_X1 U2525 ( .A1(n20197), .A2(n5363), .B1(n20205), .B2(n5080), .ZN(n2589) );
  OAI221_X1 U2526 ( .B1(n18919), .B2(n20181), .C1(n19111), .C2(n20188), .A(
        n2564), .ZN(n2562) );
  AOI22_X1 U2527 ( .A1(n20197), .A2(n5364), .B1(n20206), .B2(n5081), .ZN(n2564) );
  OAI221_X1 U2528 ( .B1(n18920), .B2(n20182), .C1(n19112), .C2(n20190), .A(
        n2539), .ZN(n2537) );
  AOI22_X1 U2529 ( .A1(n20202), .A2(n5365), .B1(n20205), .B2(n5082), .ZN(n2539) );
  OAI221_X1 U2530 ( .B1(n18921), .B2(n20182), .C1(n19113), .C2(n20189), .A(
        n2514), .ZN(n2512) );
  AOI22_X1 U2531 ( .A1(n20198), .A2(n5366), .B1(n20206), .B2(n5083), .ZN(n2514) );
  OAI221_X1 U2532 ( .B1(n18922), .B2(n20181), .C1(n19114), .C2(n20189), .A(
        n2489), .ZN(n2487) );
  AOI22_X1 U2533 ( .A1(n20198), .A2(n5367), .B1(n20206), .B2(n5084), .ZN(n2489) );
  OAI221_X1 U2534 ( .B1(n18923), .B2(n20183), .C1(n19115), .C2(n20190), .A(
        n2464), .ZN(n2462) );
  AOI22_X1 U2535 ( .A1(n20198), .A2(n5368), .B1(n20207), .B2(n5085), .ZN(n2464) );
  OAI221_X1 U2536 ( .B1(n18924), .B2(n20183), .C1(n19116), .C2(n20189), .A(
        n2439), .ZN(n2437) );
  AOI22_X1 U2537 ( .A1(n20199), .A2(n5369), .B1(n20208), .B2(n5086), .ZN(n2439) );
  OAI221_X1 U2538 ( .B1(n18925), .B2(n20185), .C1(n19117), .C2(n20192), .A(
        n2414), .ZN(n2412) );
  AOI22_X1 U2539 ( .A1(n20199), .A2(n5370), .B1(n20207), .B2(n5087), .ZN(n2414) );
  OAI221_X1 U2540 ( .B1(n18926), .B2(n20184), .C1(n19118), .C2(n20191), .A(
        n2389), .ZN(n2387) );
  AOI22_X1 U2541 ( .A1(n20200), .A2(n5371), .B1(n20208), .B2(n5088), .ZN(n2389) );
  OAI221_X1 U2542 ( .B1(n18927), .B2(n20181), .C1(n19119), .C2(n20188), .A(
        n2364), .ZN(n2362) );
  AOI22_X1 U2543 ( .A1(n20201), .A2(n5372), .B1(n20209), .B2(n5089), .ZN(n2364) );
  OAI221_X1 U2544 ( .B1(n18928), .B2(n20181), .C1(n19120), .C2(n20188), .A(
        n2339), .ZN(n2337) );
  AOI22_X1 U2545 ( .A1(n20201), .A2(n5373), .B1(n20209), .B2(n5090), .ZN(n2339) );
  OAI221_X1 U2546 ( .B1(n18929), .B2(n20182), .C1(n19121), .C2(n20189), .A(
        n2314), .ZN(n2312) );
  AOI22_X1 U2547 ( .A1(n20199), .A2(n5374), .B1(n20207), .B2(n5091), .ZN(n2314) );
  OAI221_X1 U2548 ( .B1(n18930), .B2(n20183), .C1(n19122), .C2(n20188), .A(
        n2289), .ZN(n2287) );
  AOI22_X1 U2549 ( .A1(n20200), .A2(n5375), .B1(n20208), .B2(n5092), .ZN(n2289) );
  OAI221_X1 U2550 ( .B1(n18931), .B2(n20183), .C1(n19123), .C2(n20190), .A(
        n2264), .ZN(n2262) );
  AOI22_X1 U2551 ( .A1(n20201), .A2(n5376), .B1(n20209), .B2(n5093), .ZN(n2264) );
  OAI221_X1 U2552 ( .B1(n18932), .B2(n20182), .C1(n19124), .C2(n20190), .A(
        n2239), .ZN(n2237) );
  AOI22_X1 U2553 ( .A1(n20201), .A2(n5377), .B1(n20209), .B2(n5151), .ZN(n2239) );
  OAI221_X1 U2554 ( .B1(n18933), .B2(n20186), .C1(n19125), .C2(n20191), .A(
        n2214), .ZN(n2212) );
  AOI22_X1 U2555 ( .A1(n20202), .A2(n5378), .B1(n20210), .B2(n5001), .ZN(n2214) );
  OAI221_X1 U2556 ( .B1(n18934), .B2(n20184), .C1(n19126), .C2(n20191), .A(
        n2189), .ZN(n2187) );
  AOI22_X1 U2557 ( .A1(n20202), .A2(n5379), .B1(n20210), .B2(n5002), .ZN(n2189) );
  OAI221_X1 U2558 ( .B1(n18935), .B2(n20184), .C1(n19127), .C2(n20189), .A(
        n2164), .ZN(n2162) );
  AOI22_X1 U2559 ( .A1(n20202), .A2(n5440), .B1(n20210), .B2(n5007), .ZN(n2164) );
  OAI221_X1 U2560 ( .B1(n18936), .B2(n20185), .C1(n19128), .C2(n20192), .A(
        n2139), .ZN(n2137) );
  AOI22_X1 U2561 ( .A1(n20202), .A2(n5441), .B1(n20210), .B2(n5008), .ZN(n2139) );
  OAI221_X1 U2562 ( .B1(n18937), .B2(n20184), .C1(n19129), .C2(n20193), .A(
        n2114), .ZN(n2112) );
  AOI22_X1 U2563 ( .A1(n20196), .A2(n5442), .B1(n20205), .B2(n5009), .ZN(n2114) );
  OAI221_X1 U2564 ( .B1(n18938), .B2(n20185), .C1(n19130), .C2(n20192), .A(
        n2089), .ZN(n2087) );
  AOI22_X1 U2565 ( .A1(n20196), .A2(n5443), .B1(n20209), .B2(n5010), .ZN(n2089) );
  OAI221_X1 U2566 ( .B1(n18939), .B2(n20185), .C1(n19131), .C2(n20193), .A(
        n2064), .ZN(n2062) );
  AOI22_X1 U2567 ( .A1(n20201), .A2(n5444), .B1(n20205), .B2(n5011), .ZN(n2064) );
  OAI221_X1 U2568 ( .B1(n18940), .B2(n20186), .C1(n19132), .C2(n20194), .A(
        n2039), .ZN(n2037) );
  AOI22_X1 U2569 ( .A1(n20197), .A2(n5445), .B1(n20208), .B2(n5012), .ZN(n2039) );
  OAI221_X1 U2570 ( .B1(n18941), .B2(n20186), .C1(n19133), .C2(n20194), .A(
        n2014), .ZN(n2012) );
  AOI22_X1 U2571 ( .A1(n20199), .A2(n5446), .B1(n20208), .B2(n5013), .ZN(n2014) );
  OAI221_X1 U2572 ( .B1(n18942), .B2(n20184), .C1(n19134), .C2(n20190), .A(
        n1989), .ZN(n1987) );
  AOI22_X1 U2573 ( .A1(n20196), .A2(n5447), .B1(n20210), .B2(n5014), .ZN(n1989) );
  OAI221_X1 U2574 ( .B1(n18943), .B2(n20180), .C1(n19135), .C2(n20191), .A(
        n1964), .ZN(n1962) );
  AOI22_X1 U2575 ( .A1(n20198), .A2(n5380), .B1(n20206), .B2(n5003), .ZN(n1964) );
  OAI221_X1 U2576 ( .B1(n18944), .B2(n20180), .C1(n19136), .C2(n20194), .A(
        n1939), .ZN(n1937) );
  AOI22_X1 U2577 ( .A1(n20198), .A2(n5381), .B1(n20206), .B2(n5004), .ZN(n1939) );
  OAI221_X1 U2578 ( .B1(n18945), .B2(n20185), .C1(n19137), .C2(n20193), .A(
        n1914), .ZN(n1912) );
  AOI22_X1 U2579 ( .A1(n20200), .A2(n5382), .B1(n20206), .B2(n5005), .ZN(n1914) );
  OAI221_X1 U2580 ( .B1(n18946), .B2(n20180), .C1(n19138), .C2(n20194), .A(
        n1879), .ZN(n1873) );
  AOI22_X1 U2581 ( .A1(n20200), .A2(n5383), .B1(n20207), .B2(n5006), .ZN(n1879) );
  OAI22_X1 U2582 ( .A1(n19785), .A2(n19683), .B1(n20563), .B2(n20333), .ZN(
        n3435) );
  OAI22_X1 U2583 ( .A1(n19785), .A2(n19684), .B1(n20566), .B2(n20331), .ZN(
        n3436) );
  OAI22_X1 U2584 ( .A1(n19785), .A2(n19685), .B1(n20569), .B2(n20333), .ZN(
        n3437) );
  OAI22_X1 U2585 ( .A1(n19785), .A2(n19686), .B1(n20572), .B2(n20332), .ZN(
        n3438) );
  OAI22_X1 U2586 ( .A1(n19785), .A2(n19687), .B1(n20575), .B2(n20331), .ZN(
        n3439) );
  OAI22_X1 U2587 ( .A1(n19785), .A2(n19688), .B1(n20578), .B2(n20336), .ZN(
        n3440) );
  OAI22_X1 U2588 ( .A1(n19785), .A2(n19689), .B1(n20581), .B2(n20332), .ZN(
        n3441) );
  OAI22_X1 U2589 ( .A1(n19785), .A2(n19690), .B1(n20584), .B2(n20333), .ZN(
        n3442) );
  OAI22_X1 U2590 ( .A1(n19785), .A2(n19691), .B1(n20587), .B2(n20333), .ZN(
        n3443) );
  OAI22_X1 U2591 ( .A1(n19785), .A2(n19692), .B1(n20590), .B2(n20336), .ZN(
        n3444) );
  OAI22_X1 U2592 ( .A1(n19785), .A2(n19693), .B1(n20593), .B2(n20334), .ZN(
        n3445) );
  OAI22_X1 U2593 ( .A1(n19785), .A2(n19694), .B1(n20596), .B2(n20335), .ZN(
        n3446) );
  OAI22_X1 U2594 ( .A1(n19786), .A2(n19695), .B1(n20599), .B2(n20332), .ZN(
        n3447) );
  OAI22_X1 U2595 ( .A1(n19786), .A2(n19696), .B1(n20602), .B2(n20333), .ZN(
        n3448) );
  OAI22_X1 U2596 ( .A1(n19786), .A2(n19697), .B1(n20605), .B2(n20332), .ZN(
        n3449) );
  OAI22_X1 U2597 ( .A1(n19786), .A2(n19698), .B1(n20608), .B2(n20337), .ZN(
        n3450) );
  OAI22_X1 U2598 ( .A1(n19786), .A2(n19699), .B1(n20611), .B2(n20334), .ZN(
        n3451) );
  OAI22_X1 U2599 ( .A1(n19786), .A2(n19700), .B1(n20614), .B2(n20335), .ZN(
        n3452) );
  OAI22_X1 U2600 ( .A1(n19786), .A2(n19701), .B1(n20617), .B2(n20335), .ZN(
        n3453) );
  OAI22_X1 U2601 ( .A1(n19786), .A2(n19702), .B1(n20620), .B2(n20331), .ZN(
        n3454) );
  OAI22_X1 U2602 ( .A1(n19786), .A2(n19703), .B1(n20623), .B2(n20334), .ZN(
        n3455) );
  OAI22_X1 U2603 ( .A1(n19786), .A2(n19704), .B1(n20626), .B2(n20337), .ZN(
        n3456) );
  OAI22_X1 U2604 ( .A1(n19786), .A2(n19705), .B1(n20629), .B2(n20337), .ZN(
        n3457) );
  OAI22_X1 U2605 ( .A1(n19786), .A2(n19706), .B1(n20632), .B2(n20336), .ZN(
        n3458) );
  OAI22_X1 U2606 ( .A1(n19787), .A2(n19707), .B1(n20635), .B2(n20336), .ZN(
        n3459) );
  OAI22_X1 U2607 ( .A1(n19787), .A2(n19708), .B1(n20638), .B2(n20337), .ZN(
        n3460) );
  OAI22_X1 U2608 ( .A1(n19787), .A2(n19709), .B1(n20641), .B2(n20337), .ZN(
        n3461) );
  OAI22_X1 U2609 ( .A1(n19787), .A2(n19710), .B1(n20644), .B2(n20336), .ZN(
        n3462) );
  OAI22_X1 U2610 ( .A1(n19787), .A2(n19711), .B1(n20647), .B2(n20333), .ZN(
        n3463) );
  OAI22_X1 U2611 ( .A1(n19787), .A2(n19712), .B1(n20650), .B2(n20332), .ZN(
        n3464) );
  OAI22_X1 U2612 ( .A1(n19787), .A2(n19713), .B1(n20653), .B2(n20335), .ZN(
        n3465) );
  OAI22_X1 U2613 ( .A1(n19787), .A2(n19714), .B1(n20656), .B2(n20334), .ZN(
        n3466) );
  OAI22_X1 U2614 ( .A1(n19797), .A2(n19715), .B1(n20562), .B2(n20369), .ZN(
        n3563) );
  OAI22_X1 U2615 ( .A1(n19797), .A2(n19716), .B1(n20565), .B2(n20367), .ZN(
        n3564) );
  OAI22_X1 U2616 ( .A1(n19797), .A2(n19717), .B1(n20568), .B2(n20369), .ZN(
        n3565) );
  OAI22_X1 U2617 ( .A1(n19797), .A2(n19718), .B1(n20571), .B2(n20368), .ZN(
        n3566) );
  OAI22_X1 U2618 ( .A1(n19797), .A2(n19719), .B1(n20574), .B2(n20367), .ZN(
        n3567) );
  OAI22_X1 U2619 ( .A1(n19797), .A2(n19720), .B1(n20577), .B2(n20372), .ZN(
        n3568) );
  OAI22_X1 U2620 ( .A1(n19797), .A2(n19721), .B1(n20580), .B2(n20368), .ZN(
        n3569) );
  OAI22_X1 U2621 ( .A1(n19797), .A2(n19722), .B1(n20583), .B2(n20369), .ZN(
        n3570) );
  OAI22_X1 U2622 ( .A1(n19797), .A2(n19723), .B1(n20586), .B2(n20369), .ZN(
        n3571) );
  OAI22_X1 U2623 ( .A1(n19797), .A2(n19724), .B1(n20589), .B2(n20372), .ZN(
        n3572) );
  OAI22_X1 U2624 ( .A1(n19797), .A2(n19725), .B1(n20592), .B2(n20370), .ZN(
        n3573) );
  OAI22_X1 U2625 ( .A1(n19797), .A2(n19726), .B1(n20595), .B2(n20371), .ZN(
        n3574) );
  OAI22_X1 U2626 ( .A1(n19798), .A2(n19727), .B1(n20598), .B2(n20368), .ZN(
        n3575) );
  OAI22_X1 U2627 ( .A1(n19798), .A2(n19728), .B1(n20601), .B2(n20369), .ZN(
        n3576) );
  OAI22_X1 U2628 ( .A1(n19798), .A2(n19729), .B1(n20604), .B2(n20368), .ZN(
        n3577) );
  OAI22_X1 U2629 ( .A1(n19798), .A2(n19730), .B1(n20607), .B2(n20373), .ZN(
        n3578) );
  OAI22_X1 U2630 ( .A1(n19798), .A2(n19731), .B1(n20610), .B2(n20370), .ZN(
        n3579) );
  OAI22_X1 U2631 ( .A1(n19798), .A2(n19732), .B1(n20613), .B2(n20371), .ZN(
        n3580) );
  OAI22_X1 U2632 ( .A1(n19798), .A2(n19733), .B1(n20616), .B2(n20371), .ZN(
        n3581) );
  OAI22_X1 U2633 ( .A1(n19798), .A2(n19734), .B1(n20619), .B2(n20367), .ZN(
        n3582) );
  OAI22_X1 U2634 ( .A1(n19798), .A2(n19735), .B1(n20622), .B2(n20370), .ZN(
        n3583) );
  OAI22_X1 U2635 ( .A1(n19798), .A2(n19736), .B1(n20625), .B2(n20373), .ZN(
        n3584) );
  OAI22_X1 U2636 ( .A1(n19798), .A2(n19737), .B1(n20628), .B2(n20373), .ZN(
        n3585) );
  OAI22_X1 U2637 ( .A1(n19798), .A2(n19738), .B1(n20631), .B2(n20372), .ZN(
        n3586) );
  OAI22_X1 U2638 ( .A1(n19799), .A2(n19739), .B1(n20634), .B2(n20372), .ZN(
        n3587) );
  OAI22_X1 U2639 ( .A1(n19799), .A2(n19740), .B1(n20637), .B2(n20373), .ZN(
        n3588) );
  OAI22_X1 U2640 ( .A1(n19799), .A2(n19741), .B1(n20640), .B2(n20373), .ZN(
        n3589) );
  OAI22_X1 U2641 ( .A1(n19799), .A2(n19742), .B1(n20643), .B2(n20372), .ZN(
        n3590) );
  OAI22_X1 U2642 ( .A1(n19799), .A2(n19743), .B1(n20646), .B2(n20369), .ZN(
        n3591) );
  OAI22_X1 U2643 ( .A1(n19799), .A2(n19744), .B1(n20649), .B2(n20368), .ZN(
        n3592) );
  OAI22_X1 U2644 ( .A1(n19799), .A2(n19745), .B1(n20652), .B2(n20371), .ZN(
        n3593) );
  OAI22_X1 U2645 ( .A1(n19799), .A2(n19746), .B1(n20655), .B2(n20370), .ZN(
        n3594) );
  OAI22_X1 U2646 ( .A1(n5479), .A2(n19800), .B1(n20562), .B2(n20376), .ZN(
        n3595) );
  OAI22_X1 U2647 ( .A1(n5480), .A2(n19800), .B1(n20565), .B2(n20375), .ZN(
        n3596) );
  OAI22_X1 U2648 ( .A1(n5481), .A2(n19800), .B1(n20568), .B2(n20376), .ZN(
        n3597) );
  OAI22_X1 U2649 ( .A1(n5482), .A2(n19800), .B1(n20571), .B2(n20378), .ZN(
        n3598) );
  OAI22_X1 U2650 ( .A1(n5483), .A2(n19800), .B1(n20574), .B2(n20376), .ZN(
        n3599) );
  OAI22_X1 U2651 ( .A1(n5484), .A2(n19800), .B1(n20577), .B2(n20381), .ZN(
        n3600) );
  OAI22_X1 U2652 ( .A1(n5485), .A2(n19800), .B1(n20580), .B2(n20377), .ZN(
        n3601) );
  OAI22_X1 U2653 ( .A1(n5486), .A2(n19800), .B1(n20583), .B2(n20378), .ZN(
        n3602) );
  OAI22_X1 U2654 ( .A1(n5487), .A2(n19800), .B1(n20586), .B2(n20378), .ZN(
        n3603) );
  OAI22_X1 U2655 ( .A1(n5488), .A2(n19800), .B1(n20589), .B2(n20380), .ZN(
        n3604) );
  OAI22_X1 U2656 ( .A1(n5489), .A2(n19800), .B1(n20592), .B2(n20379), .ZN(
        n3605) );
  OAI22_X1 U2657 ( .A1(n5490), .A2(n19800), .B1(n20595), .B2(n20380), .ZN(
        n3606) );
  OAI22_X1 U2658 ( .A1(n5491), .A2(n19801), .B1(n20598), .B2(n20377), .ZN(
        n3607) );
  OAI22_X1 U2659 ( .A1(n5492), .A2(n19801), .B1(n20601), .B2(n20378), .ZN(
        n3608) );
  OAI22_X1 U2660 ( .A1(n5493), .A2(n19801), .B1(n20604), .B2(n20377), .ZN(
        n3609) );
  OAI22_X1 U2661 ( .A1(n5494), .A2(n19801), .B1(n20607), .B2(n20379), .ZN(
        n3610) );
  OAI22_X1 U2662 ( .A1(n5495), .A2(n19801), .B1(n20610), .B2(n20379), .ZN(
        n3611) );
  OAI22_X1 U2663 ( .A1(n5496), .A2(n19801), .B1(n20613), .B2(n20380), .ZN(
        n3612) );
  OAI22_X1 U2664 ( .A1(n5497), .A2(n19801), .B1(n20616), .B2(n20380), .ZN(
        n3613) );
  OAI22_X1 U2665 ( .A1(n5498), .A2(n19801), .B1(n20619), .B2(n20376), .ZN(
        n3614) );
  OAI22_X1 U2666 ( .A1(n5499), .A2(n19801), .B1(n20622), .B2(n20379), .ZN(
        n3615) );
  OAI22_X1 U2667 ( .A1(n5500), .A2(n19801), .B1(n20625), .B2(n20382), .ZN(
        n3616) );
  OAI22_X1 U2668 ( .A1(n5501), .A2(n19801), .B1(n20628), .B2(n20382), .ZN(
        n3617) );
  OAI22_X1 U2669 ( .A1(n5475), .A2(n19801), .B1(n20631), .B2(n20381), .ZN(
        n3618) );
  OAI22_X1 U2670 ( .A1(n5502), .A2(n19802), .B1(n20634), .B2(n20381), .ZN(
        n3619) );
  OAI22_X1 U2671 ( .A1(n5503), .A2(n19802), .B1(n20637), .B2(n20382), .ZN(
        n3620) );
  OAI22_X1 U2672 ( .A1(n5504), .A2(n19802), .B1(n20640), .B2(n20382), .ZN(
        n3621) );
  OAI22_X1 U2673 ( .A1(n5505), .A2(n19802), .B1(n20643), .B2(n20381), .ZN(
        n3622) );
  OAI22_X1 U2674 ( .A1(n5506), .A2(n19802), .B1(n20646), .B2(n20375), .ZN(
        n3623) );
  OAI22_X1 U2675 ( .A1(n5507), .A2(n19802), .B1(n20649), .B2(n20375), .ZN(
        n3624) );
  OAI22_X1 U2676 ( .A1(n5508), .A2(n19802), .B1(n20652), .B2(n20375), .ZN(
        n3625) );
  OAI22_X1 U2677 ( .A1(n5509), .A2(n19802), .B1(n20655), .B2(n20377), .ZN(
        n3626) );
  OAI22_X1 U2678 ( .A1(n19803), .A2(n19651), .B1(n20562), .B2(n20387), .ZN(
        n3627) );
  OAI22_X1 U2679 ( .A1(n19803), .A2(n19652), .B1(n20565), .B2(n20385), .ZN(
        n3628) );
  OAI22_X1 U2680 ( .A1(n19803), .A2(n19653), .B1(n20568), .B2(n20387), .ZN(
        n3629) );
  OAI22_X1 U2681 ( .A1(n19803), .A2(n19654), .B1(n20571), .B2(n20386), .ZN(
        n3630) );
  OAI22_X1 U2682 ( .A1(n19803), .A2(n19655), .B1(n20574), .B2(n20385), .ZN(
        n3631) );
  OAI22_X1 U2683 ( .A1(n19803), .A2(n19656), .B1(n20577), .B2(n20390), .ZN(
        n3632) );
  OAI22_X1 U2684 ( .A1(n19803), .A2(n19657), .B1(n20580), .B2(n20386), .ZN(
        n3633) );
  OAI22_X1 U2685 ( .A1(n19803), .A2(n19658), .B1(n20583), .B2(n20387), .ZN(
        n3634) );
  OAI22_X1 U2686 ( .A1(n19803), .A2(n19659), .B1(n20586), .B2(n20387), .ZN(
        n3635) );
  OAI22_X1 U2687 ( .A1(n19803), .A2(n19660), .B1(n20589), .B2(n20390), .ZN(
        n3636) );
  OAI22_X1 U2688 ( .A1(n19803), .A2(n19661), .B1(n20592), .B2(n20388), .ZN(
        n3637) );
  OAI22_X1 U2689 ( .A1(n19803), .A2(n19662), .B1(n20595), .B2(n20389), .ZN(
        n3638) );
  OAI22_X1 U2690 ( .A1(n19804), .A2(n19663), .B1(n20598), .B2(n20386), .ZN(
        n3639) );
  OAI22_X1 U2691 ( .A1(n19804), .A2(n19664), .B1(n20601), .B2(n20387), .ZN(
        n3640) );
  OAI22_X1 U2692 ( .A1(n19804), .A2(n19665), .B1(n20604), .B2(n20386), .ZN(
        n3641) );
  OAI22_X1 U2693 ( .A1(n19804), .A2(n19666), .B1(n20607), .B2(n20391), .ZN(
        n3642) );
  OAI22_X1 U2694 ( .A1(n19804), .A2(n19667), .B1(n20610), .B2(n20388), .ZN(
        n3643) );
  OAI22_X1 U2695 ( .A1(n19804), .A2(n19668), .B1(n20613), .B2(n20389), .ZN(
        n3644) );
  OAI22_X1 U2696 ( .A1(n19804), .A2(n19669), .B1(n20616), .B2(n20389), .ZN(
        n3645) );
  OAI22_X1 U2697 ( .A1(n19804), .A2(n19670), .B1(n20619), .B2(n20385), .ZN(
        n3646) );
  OAI22_X1 U2698 ( .A1(n19804), .A2(n19671), .B1(n20622), .B2(n20388), .ZN(
        n3647) );
  OAI22_X1 U2699 ( .A1(n19804), .A2(n19672), .B1(n20625), .B2(n20391), .ZN(
        n3648) );
  OAI22_X1 U2700 ( .A1(n19804), .A2(n19673), .B1(n20628), .B2(n20391), .ZN(
        n3649) );
  OAI22_X1 U2701 ( .A1(n19804), .A2(n19674), .B1(n20631), .B2(n20390), .ZN(
        n3650) );
  OAI22_X1 U2702 ( .A1(n19805), .A2(n19675), .B1(n20634), .B2(n20390), .ZN(
        n3651) );
  OAI22_X1 U2703 ( .A1(n19805), .A2(n19676), .B1(n20637), .B2(n20391), .ZN(
        n3652) );
  OAI22_X1 U2704 ( .A1(n19805), .A2(n19677), .B1(n20640), .B2(n20391), .ZN(
        n3653) );
  OAI22_X1 U2705 ( .A1(n19805), .A2(n19678), .B1(n20643), .B2(n20390), .ZN(
        n3654) );
  OAI22_X1 U2706 ( .A1(n19805), .A2(n19679), .B1(n20646), .B2(n20387), .ZN(
        n3655) );
  OAI22_X1 U2707 ( .A1(n19805), .A2(n19680), .B1(n20649), .B2(n20386), .ZN(
        n3656) );
  OAI22_X1 U2708 ( .A1(n19805), .A2(n19681), .B1(n20652), .B2(n20389), .ZN(
        n3657) );
  OAI22_X1 U2709 ( .A1(n19805), .A2(n19682), .B1(n20655), .B2(n20388), .ZN(
        n3658) );
  OAI22_X1 U2710 ( .A1(n8486), .A2(n19815), .B1(n20562), .B2(n20421), .ZN(
        n3755) );
  OAI22_X1 U2711 ( .A1(n8487), .A2(n19815), .B1(n20565), .B2(n20420), .ZN(
        n3756) );
  OAI22_X1 U2712 ( .A1(n8488), .A2(n19815), .B1(n20568), .B2(n20421), .ZN(
        n3757) );
  OAI22_X1 U2713 ( .A1(n8489), .A2(n19815), .B1(n20571), .B2(n20423), .ZN(
        n3758) );
  OAI22_X1 U2714 ( .A1(n8490), .A2(n19815), .B1(n20574), .B2(n20421), .ZN(
        n3759) );
  OAI22_X1 U2715 ( .A1(n8491), .A2(n19815), .B1(n20577), .B2(n20426), .ZN(
        n3760) );
  OAI22_X1 U2716 ( .A1(n8492), .A2(n19815), .B1(n20580), .B2(n20422), .ZN(
        n3761) );
  OAI22_X1 U2717 ( .A1(n8493), .A2(n19815), .B1(n20583), .B2(n20423), .ZN(
        n3762) );
  OAI22_X1 U2718 ( .A1(n8494), .A2(n19815), .B1(n20586), .B2(n20423), .ZN(
        n3763) );
  OAI22_X1 U2719 ( .A1(n8495), .A2(n19815), .B1(n20589), .B2(n20425), .ZN(
        n3764) );
  OAI22_X1 U2720 ( .A1(n8496), .A2(n19815), .B1(n20592), .B2(n20424), .ZN(
        n3765) );
  OAI22_X1 U2721 ( .A1(n8497), .A2(n19815), .B1(n20595), .B2(n20425), .ZN(
        n3766) );
  OAI22_X1 U2722 ( .A1(n8498), .A2(n19816), .B1(n20598), .B2(n20422), .ZN(
        n3767) );
  OAI22_X1 U2723 ( .A1(n8499), .A2(n19816), .B1(n20601), .B2(n20423), .ZN(
        n3768) );
  OAI22_X1 U2724 ( .A1(n8500), .A2(n19816), .B1(n20604), .B2(n20422), .ZN(
        n3769) );
  OAI22_X1 U2725 ( .A1(n8501), .A2(n19816), .B1(n20607), .B2(n20424), .ZN(
        n3770) );
  OAI22_X1 U2726 ( .A1(n8502), .A2(n19816), .B1(n20610), .B2(n20424), .ZN(
        n3771) );
  OAI22_X1 U2727 ( .A1(n8503), .A2(n19816), .B1(n20613), .B2(n20425), .ZN(
        n3772) );
  OAI22_X1 U2728 ( .A1(n8504), .A2(n19816), .B1(n20616), .B2(n20425), .ZN(
        n3773) );
  OAI22_X1 U2729 ( .A1(n8505), .A2(n19816), .B1(n20619), .B2(n20421), .ZN(
        n3774) );
  OAI22_X1 U2730 ( .A1(n8506), .A2(n19816), .B1(n20622), .B2(n20424), .ZN(
        n3775) );
  OAI22_X1 U2731 ( .A1(n8507), .A2(n19816), .B1(n20625), .B2(n20427), .ZN(
        n3776) );
  OAI22_X1 U2732 ( .A1(n8508), .A2(n19816), .B1(n20628), .B2(n20427), .ZN(
        n3777) );
  OAI22_X1 U2733 ( .A1(n8509), .A2(n19816), .B1(n20631), .B2(n20426), .ZN(
        n3778) );
  OAI22_X1 U2734 ( .A1(n8510), .A2(n19817), .B1(n20634), .B2(n20426), .ZN(
        n3779) );
  OAI22_X1 U2735 ( .A1(n8511), .A2(n19817), .B1(n20637), .B2(n20427), .ZN(
        n3780) );
  OAI22_X1 U2736 ( .A1(n8512), .A2(n19817), .B1(n20640), .B2(n20427), .ZN(
        n3781) );
  OAI22_X1 U2737 ( .A1(n8513), .A2(n19817), .B1(n20643), .B2(n20426), .ZN(
        n3782) );
  OAI22_X1 U2738 ( .A1(n8514), .A2(n19817), .B1(n20646), .B2(n20420), .ZN(
        n3783) );
  OAI22_X1 U2739 ( .A1(n8515), .A2(n19817), .B1(n20649), .B2(n20420), .ZN(
        n3784) );
  OAI22_X1 U2740 ( .A1(n8516), .A2(n19817), .B1(n20652), .B2(n20420), .ZN(
        n3785) );
  OAI22_X1 U2741 ( .A1(n8517), .A2(n19817), .B1(n20655), .B2(n20422), .ZN(
        n3786) );
  OAI22_X1 U2742 ( .A1(n5510), .A2(n19824), .B1(n20562), .B2(n20448), .ZN(
        n3851) );
  OAI22_X1 U2743 ( .A1(n5511), .A2(n19824), .B1(n20565), .B2(n20447), .ZN(
        n3852) );
  OAI22_X1 U2744 ( .A1(n5512), .A2(n19824), .B1(n20568), .B2(n20448), .ZN(
        n3853) );
  OAI22_X1 U2745 ( .A1(n5513), .A2(n19824), .B1(n20571), .B2(n20450), .ZN(
        n3854) );
  OAI22_X1 U2746 ( .A1(n5514), .A2(n19824), .B1(n20574), .B2(n20448), .ZN(
        n3855) );
  OAI22_X1 U2747 ( .A1(n5515), .A2(n19824), .B1(n20577), .B2(n20453), .ZN(
        n3856) );
  OAI22_X1 U2748 ( .A1(n5516), .A2(n19824), .B1(n20580), .B2(n20449), .ZN(
        n3857) );
  OAI22_X1 U2749 ( .A1(n5517), .A2(n19824), .B1(n20583), .B2(n20450), .ZN(
        n3858) );
  OAI22_X1 U2750 ( .A1(n5518), .A2(n19824), .B1(n20586), .B2(n20450), .ZN(
        n3859) );
  OAI22_X1 U2751 ( .A1(n5519), .A2(n19824), .B1(n20589), .B2(n20452), .ZN(
        n3860) );
  OAI22_X1 U2752 ( .A1(n5520), .A2(n19824), .B1(n20592), .B2(n20451), .ZN(
        n3861) );
  OAI22_X1 U2753 ( .A1(n5521), .A2(n19824), .B1(n20595), .B2(n20452), .ZN(
        n3862) );
  OAI22_X1 U2754 ( .A1(n5522), .A2(n19825), .B1(n20598), .B2(n20449), .ZN(
        n3863) );
  OAI22_X1 U2755 ( .A1(n5523), .A2(n19825), .B1(n20601), .B2(n20450), .ZN(
        n3864) );
  OAI22_X1 U2756 ( .A1(n5524), .A2(n19825), .B1(n20604), .B2(n20449), .ZN(
        n3865) );
  OAI22_X1 U2757 ( .A1(n5525), .A2(n19825), .B1(n20607), .B2(n20451), .ZN(
        n3866) );
  OAI22_X1 U2758 ( .A1(n5526), .A2(n19825), .B1(n20610), .B2(n20451), .ZN(
        n3867) );
  OAI22_X1 U2759 ( .A1(n5527), .A2(n19825), .B1(n20613), .B2(n20452), .ZN(
        n3868) );
  OAI22_X1 U2760 ( .A1(n5528), .A2(n19825), .B1(n20616), .B2(n20452), .ZN(
        n3869) );
  OAI22_X1 U2761 ( .A1(n5529), .A2(n19825), .B1(n20619), .B2(n20448), .ZN(
        n3870) );
  OAI22_X1 U2762 ( .A1(n5530), .A2(n19825), .B1(n20622), .B2(n20451), .ZN(
        n3871) );
  OAI22_X1 U2763 ( .A1(n5531), .A2(n19825), .B1(n20625), .B2(n20454), .ZN(
        n3872) );
  OAI22_X1 U2764 ( .A1(n5532), .A2(n19825), .B1(n20628), .B2(n20454), .ZN(
        n3873) );
  OAI22_X1 U2765 ( .A1(n5476), .A2(n19825), .B1(n20631), .B2(n20453), .ZN(
        n3874) );
  OAI22_X1 U2766 ( .A1(n5533), .A2(n19826), .B1(n20634), .B2(n20453), .ZN(
        n3875) );
  OAI22_X1 U2767 ( .A1(n5534), .A2(n19826), .B1(n20637), .B2(n20454), .ZN(
        n3876) );
  OAI22_X1 U2768 ( .A1(n5535), .A2(n19826), .B1(n20640), .B2(n20454), .ZN(
        n3877) );
  OAI22_X1 U2769 ( .A1(n5536), .A2(n19826), .B1(n20643), .B2(n20453), .ZN(
        n3878) );
  OAI22_X1 U2770 ( .A1(n5537), .A2(n19826), .B1(n20646), .B2(n20447), .ZN(
        n3879) );
  OAI22_X1 U2771 ( .A1(n5538), .A2(n19826), .B1(n20649), .B2(n20447), .ZN(
        n3880) );
  OAI22_X1 U2772 ( .A1(n5539), .A2(n19826), .B1(n20652), .B2(n20447), .ZN(
        n3881) );
  OAI22_X1 U2773 ( .A1(n5540), .A2(n19826), .B1(n20655), .B2(n20449), .ZN(
        n3882) );
  OAI22_X1 U2774 ( .A1(n4952), .A2(n19827), .B1(n20562), .B2(n20457), .ZN(
        n3883) );
  OAI22_X1 U2775 ( .A1(n4953), .A2(n19827), .B1(n20565), .B2(n20456), .ZN(
        n3884) );
  OAI22_X1 U2776 ( .A1(n4954), .A2(n19827), .B1(n20568), .B2(n20457), .ZN(
        n3885) );
  OAI22_X1 U2777 ( .A1(n4955), .A2(n19827), .B1(n20571), .B2(n20459), .ZN(
        n3886) );
  OAI22_X1 U2778 ( .A1(n4956), .A2(n19827), .B1(n20574), .B2(n20457), .ZN(
        n3887) );
  OAI22_X1 U2779 ( .A1(n4957), .A2(n19827), .B1(n20577), .B2(n20462), .ZN(
        n3888) );
  OAI22_X1 U2780 ( .A1(n4958), .A2(n19827), .B1(n20580), .B2(n20458), .ZN(
        n3889) );
  OAI22_X1 U2781 ( .A1(n4959), .A2(n19827), .B1(n20583), .B2(n20459), .ZN(
        n3890) );
  OAI22_X1 U2782 ( .A1(n4960), .A2(n19827), .B1(n20586), .B2(n20459), .ZN(
        n3891) );
  OAI22_X1 U2783 ( .A1(n4961), .A2(n19827), .B1(n20589), .B2(n20461), .ZN(
        n3892) );
  OAI22_X1 U2784 ( .A1(n4962), .A2(n19827), .B1(n20592), .B2(n20460), .ZN(
        n3893) );
  OAI22_X1 U2785 ( .A1(n4963), .A2(n19827), .B1(n20595), .B2(n20461), .ZN(
        n3894) );
  OAI22_X1 U2786 ( .A1(n4964), .A2(n19828), .B1(n20598), .B2(n20458), .ZN(
        n3895) );
  OAI22_X1 U2787 ( .A1(n4965), .A2(n19828), .B1(n20601), .B2(n20459), .ZN(
        n3896) );
  OAI22_X1 U2788 ( .A1(n4966), .A2(n19828), .B1(n20604), .B2(n20458), .ZN(
        n3897) );
  OAI22_X1 U2789 ( .A1(n4967), .A2(n19828), .B1(n20607), .B2(n20460), .ZN(
        n3898) );
  OAI22_X1 U2790 ( .A1(n4968), .A2(n19828), .B1(n20610), .B2(n20460), .ZN(
        n3899) );
  OAI22_X1 U2791 ( .A1(n4969), .A2(n19828), .B1(n20613), .B2(n20461), .ZN(
        n3900) );
  OAI22_X1 U2792 ( .A1(n4970), .A2(n19828), .B1(n20616), .B2(n20461), .ZN(
        n3901) );
  OAI22_X1 U2793 ( .A1(n4971), .A2(n19828), .B1(n20619), .B2(n20457), .ZN(
        n3902) );
  OAI22_X1 U2794 ( .A1(n4972), .A2(n19828), .B1(n20622), .B2(n20460), .ZN(
        n3903) );
  OAI22_X1 U2795 ( .A1(n4973), .A2(n19828), .B1(n20625), .B2(n20463), .ZN(
        n3904) );
  OAI22_X1 U2796 ( .A1(n4974), .A2(n19828), .B1(n20628), .B2(n20463), .ZN(
        n3905) );
  OAI22_X1 U2797 ( .A1(n4975), .A2(n19828), .B1(n20631), .B2(n20462), .ZN(
        n3906) );
  OAI22_X1 U2798 ( .A1(n4977), .A2(n19829), .B1(n20634), .B2(n20462), .ZN(
        n3907) );
  OAI22_X1 U2799 ( .A1(n4882), .A2(n19829), .B1(n20637), .B2(n20463), .ZN(
        n3908) );
  OAI22_X1 U2800 ( .A1(n4883), .A2(n19829), .B1(n20640), .B2(n20463), .ZN(
        n3909) );
  OAI22_X1 U2801 ( .A1(n4884), .A2(n19829), .B1(n20643), .B2(n20462), .ZN(
        n3910) );
  OAI22_X1 U2802 ( .A1(n4885), .A2(n19829), .B1(n20646), .B2(n20456), .ZN(
        n3911) );
  OAI22_X1 U2803 ( .A1(n4886), .A2(n19829), .B1(n20649), .B2(n20456), .ZN(
        n3912) );
  OAI22_X1 U2804 ( .A1(n4887), .A2(n19829), .B1(n20652), .B2(n20456), .ZN(
        n3913) );
  OAI22_X1 U2805 ( .A1(n4888), .A2(n19829), .B1(n20655), .B2(n20458), .ZN(
        n3914) );
  OAI22_X1 U2806 ( .A1(n5541), .A2(n19830), .B1(n20562), .B2(n20466), .ZN(
        n3915) );
  OAI22_X1 U2807 ( .A1(n5542), .A2(n19830), .B1(n20565), .B2(n20465), .ZN(
        n3916) );
  OAI22_X1 U2808 ( .A1(n5543), .A2(n19830), .B1(n20568), .B2(n20466), .ZN(
        n3917) );
  OAI22_X1 U2809 ( .A1(n5544), .A2(n19830), .B1(n20571), .B2(n20468), .ZN(
        n3918) );
  OAI22_X1 U2810 ( .A1(n5545), .A2(n19830), .B1(n20574), .B2(n20466), .ZN(
        n3919) );
  OAI22_X1 U2811 ( .A1(n5546), .A2(n19830), .B1(n20577), .B2(n20471), .ZN(
        n3920) );
  OAI22_X1 U2812 ( .A1(n5547), .A2(n19830), .B1(n20580), .B2(n20467), .ZN(
        n3921) );
  OAI22_X1 U2813 ( .A1(n5548), .A2(n19830), .B1(n20583), .B2(n20468), .ZN(
        n3922) );
  OAI22_X1 U2814 ( .A1(n5549), .A2(n19830), .B1(n20586), .B2(n20468), .ZN(
        n3923) );
  OAI22_X1 U2815 ( .A1(n5550), .A2(n19830), .B1(n20589), .B2(n20470), .ZN(
        n3924) );
  OAI22_X1 U2816 ( .A1(n5551), .A2(n19830), .B1(n20592), .B2(n20469), .ZN(
        n3925) );
  OAI22_X1 U2817 ( .A1(n5552), .A2(n19830), .B1(n20595), .B2(n20470), .ZN(
        n3926) );
  OAI22_X1 U2818 ( .A1(n5553), .A2(n19831), .B1(n20598), .B2(n20467), .ZN(
        n3927) );
  OAI22_X1 U2819 ( .A1(n5554), .A2(n19831), .B1(n20601), .B2(n20468), .ZN(
        n3928) );
  OAI22_X1 U2820 ( .A1(n5555), .A2(n19831), .B1(n20604), .B2(n20467), .ZN(
        n3929) );
  OAI22_X1 U2821 ( .A1(n5556), .A2(n19831), .B1(n20607), .B2(n20469), .ZN(
        n3930) );
  OAI22_X1 U2822 ( .A1(n5557), .A2(n19831), .B1(n20610), .B2(n20469), .ZN(
        n3931) );
  OAI22_X1 U2823 ( .A1(n5558), .A2(n19831), .B1(n20613), .B2(n20470), .ZN(
        n3932) );
  OAI22_X1 U2824 ( .A1(n5559), .A2(n19831), .B1(n20616), .B2(n20470), .ZN(
        n3933) );
  OAI22_X1 U2825 ( .A1(n5560), .A2(n19831), .B1(n20619), .B2(n20466), .ZN(
        n3934) );
  OAI22_X1 U2826 ( .A1(n5561), .A2(n19831), .B1(n20622), .B2(n20469), .ZN(
        n3935) );
  OAI22_X1 U2827 ( .A1(n5562), .A2(n19831), .B1(n20625), .B2(n20472), .ZN(
        n3936) );
  OAI22_X1 U2828 ( .A1(n5563), .A2(n19831), .B1(n20628), .B2(n20472), .ZN(
        n3937) );
  OAI22_X1 U2829 ( .A1(n5477), .A2(n19831), .B1(n20631), .B2(n20471), .ZN(
        n3938) );
  OAI22_X1 U2830 ( .A1(n5564), .A2(n19832), .B1(n20634), .B2(n20471), .ZN(
        n3939) );
  OAI22_X1 U2831 ( .A1(n5565), .A2(n19832), .B1(n20637), .B2(n20472), .ZN(
        n3940) );
  OAI22_X1 U2832 ( .A1(n5566), .A2(n19832), .B1(n20640), .B2(n20472), .ZN(
        n3941) );
  OAI22_X1 U2833 ( .A1(n5567), .A2(n19832), .B1(n20643), .B2(n20471), .ZN(
        n3942) );
  OAI22_X1 U2834 ( .A1(n5568), .A2(n19832), .B1(n20646), .B2(n20465), .ZN(
        n3943) );
  OAI22_X1 U2835 ( .A1(n5569), .A2(n19832), .B1(n20649), .B2(n20465), .ZN(
        n3944) );
  OAI22_X1 U2836 ( .A1(n5570), .A2(n19832), .B1(n20652), .B2(n20465), .ZN(
        n3945) );
  OAI22_X1 U2837 ( .A1(n5571), .A2(n19832), .B1(n20655), .B2(n20467), .ZN(
        n3946) );
  OAI22_X1 U2838 ( .A1(n5572), .A2(n19839), .B1(n20561), .B2(n20490), .ZN(
        n4011) );
  OAI22_X1 U2839 ( .A1(n5573), .A2(n19839), .B1(n20564), .B2(n20491), .ZN(
        n4012) );
  OAI22_X1 U2840 ( .A1(n5574), .A2(n19839), .B1(n20567), .B2(n20490), .ZN(
        n4013) );
  OAI22_X1 U2841 ( .A1(n5575), .A2(n19839), .B1(n20570), .B2(n20491), .ZN(
        n4014) );
  OAI22_X1 U2842 ( .A1(n5576), .A2(n19839), .B1(n20573), .B2(n20492), .ZN(
        n4015) );
  OAI22_X1 U2843 ( .A1(n5577), .A2(n19839), .B1(n20576), .B2(n20490), .ZN(
        n4016) );
  OAI22_X1 U2844 ( .A1(n5578), .A2(n19839), .B1(n20579), .B2(n20492), .ZN(
        n4017) );
  OAI22_X1 U2845 ( .A1(n5579), .A2(n19839), .B1(n20582), .B2(n20493), .ZN(
        n4018) );
  OAI22_X1 U2846 ( .A1(n5580), .A2(n19839), .B1(n20585), .B2(n20493), .ZN(
        n4019) );
  OAI22_X1 U2847 ( .A1(n5581), .A2(n19839), .B1(n20588), .B2(n20494), .ZN(
        n4020) );
  OAI22_X1 U2848 ( .A1(n5582), .A2(n19839), .B1(n20591), .B2(n20495), .ZN(
        n4021) );
  OAI22_X1 U2849 ( .A1(n5583), .A2(n19839), .B1(n20594), .B2(n20491), .ZN(
        n4022) );
  OAI22_X1 U2850 ( .A1(n5584), .A2(n19840), .B1(n20597), .B2(n20494), .ZN(
        n4023) );
  OAI22_X1 U2851 ( .A1(n5585), .A2(n19840), .B1(n20600), .B2(n20495), .ZN(
        n4024) );
  OAI22_X1 U2852 ( .A1(n5586), .A2(n19840), .B1(n20603), .B2(n20490), .ZN(
        n4025) );
  OAI22_X1 U2853 ( .A1(n5587), .A2(n19840), .B1(n20606), .B2(n20491), .ZN(
        n4026) );
  OAI22_X1 U2854 ( .A1(n5588), .A2(n19840), .B1(n20609), .B2(n20492), .ZN(
        n4027) );
  OAI22_X1 U2855 ( .A1(n5589), .A2(n19840), .B1(n20612), .B2(n20492), .ZN(
        n4028) );
  OAI22_X1 U2856 ( .A1(n5590), .A2(n19840), .B1(n20615), .B2(n20490), .ZN(
        n4029) );
  OAI22_X1 U2857 ( .A1(n5591), .A2(n19840), .B1(n20618), .B2(n20491), .ZN(
        n4030) );
  OAI22_X1 U2858 ( .A1(n5592), .A2(n19840), .B1(n20621), .B2(n20493), .ZN(
        n4031) );
  OAI22_X1 U2859 ( .A1(n5593), .A2(n19840), .B1(n20624), .B2(n20494), .ZN(
        n4032) );
  OAI22_X1 U2860 ( .A1(n5594), .A2(n19840), .B1(n20627), .B2(n20495), .ZN(
        n4033) );
  OAI22_X1 U2861 ( .A1(n5478), .A2(n19840), .B1(n20630), .B2(n20493), .ZN(
        n4034) );
  OAI22_X1 U2862 ( .A1(n5595), .A2(n19841), .B1(n20633), .B2(n20492), .ZN(
        n4035) );
  OAI22_X1 U2863 ( .A1(n5596), .A2(n19841), .B1(n20636), .B2(n20493), .ZN(
        n4036) );
  OAI22_X1 U2864 ( .A1(n5597), .A2(n19841), .B1(n20639), .B2(n20490), .ZN(
        n4037) );
  OAI22_X1 U2865 ( .A1(n5598), .A2(n19841), .B1(n20642), .B2(n20491), .ZN(
        n4038) );
  OAI22_X1 U2866 ( .A1(n5599), .A2(n19841), .B1(n20645), .B2(n20492), .ZN(
        n4039) );
  OAI22_X1 U2867 ( .A1(n5600), .A2(n19841), .B1(n20648), .B2(n20494), .ZN(
        n4040) );
  OAI22_X1 U2868 ( .A1(n5601), .A2(n19841), .B1(n20651), .B2(n20494), .ZN(
        n4041) );
  OAI22_X1 U2869 ( .A1(n5602), .A2(n19841), .B1(n20654), .B2(n20495), .ZN(
        n4042) );
  OAI22_X1 U2870 ( .A1(n19842), .A2(n19747), .B1(n20561), .B2(n20500), .ZN(
        n4043) );
  OAI22_X1 U2871 ( .A1(n19842), .A2(n19748), .B1(n20564), .B2(n20498), .ZN(
        n4044) );
  OAI22_X1 U2872 ( .A1(n19842), .A2(n19749), .B1(n20567), .B2(n20500), .ZN(
        n4045) );
  OAI22_X1 U2873 ( .A1(n19842), .A2(n19750), .B1(n20570), .B2(n20499), .ZN(
        n4046) );
  OAI22_X1 U2874 ( .A1(n19842), .A2(n19751), .B1(n20573), .B2(n20498), .ZN(
        n4047) );
  OAI22_X1 U2875 ( .A1(n19842), .A2(n19752), .B1(n20576), .B2(n20503), .ZN(
        n4048) );
  OAI22_X1 U2876 ( .A1(n19842), .A2(n19753), .B1(n20579), .B2(n20499), .ZN(
        n4049) );
  OAI22_X1 U2877 ( .A1(n19842), .A2(n19754), .B1(n20582), .B2(n20500), .ZN(
        n4050) );
  OAI22_X1 U2878 ( .A1(n19842), .A2(n19755), .B1(n20585), .B2(n20500), .ZN(
        n4051) );
  OAI22_X1 U2879 ( .A1(n19842), .A2(n19756), .B1(n20588), .B2(n20503), .ZN(
        n4052) );
  OAI22_X1 U2880 ( .A1(n19842), .A2(n19757), .B1(n20591), .B2(n20501), .ZN(
        n4053) );
  OAI22_X1 U2881 ( .A1(n19842), .A2(n19758), .B1(n20594), .B2(n20502), .ZN(
        n4054) );
  OAI22_X1 U2882 ( .A1(n19843), .A2(n19759), .B1(n20597), .B2(n20499), .ZN(
        n4055) );
  OAI22_X1 U2883 ( .A1(n19843), .A2(n19760), .B1(n20600), .B2(n20500), .ZN(
        n4056) );
  OAI22_X1 U2884 ( .A1(n19843), .A2(n19761), .B1(n20603), .B2(n20499), .ZN(
        n4057) );
  OAI22_X1 U2885 ( .A1(n19843), .A2(n19762), .B1(n20606), .B2(n20504), .ZN(
        n4058) );
  OAI22_X1 U2886 ( .A1(n19843), .A2(n19763), .B1(n20609), .B2(n20501), .ZN(
        n4059) );
  OAI22_X1 U2887 ( .A1(n19843), .A2(n19764), .B1(n20612), .B2(n20502), .ZN(
        n4060) );
  OAI22_X1 U2888 ( .A1(n19843), .A2(n19765), .B1(n20615), .B2(n20502), .ZN(
        n4061) );
  OAI22_X1 U2889 ( .A1(n19843), .A2(n19766), .B1(n20618), .B2(n20498), .ZN(
        n4062) );
  OAI22_X1 U2890 ( .A1(n19843), .A2(n19767), .B1(n20621), .B2(n20501), .ZN(
        n4063) );
  OAI22_X1 U2891 ( .A1(n19843), .A2(n19768), .B1(n20624), .B2(n20504), .ZN(
        n4064) );
  OAI22_X1 U2892 ( .A1(n19843), .A2(n19769), .B1(n20627), .B2(n20504), .ZN(
        n4065) );
  OAI22_X1 U2893 ( .A1(n19843), .A2(n19770), .B1(n20630), .B2(n20503), .ZN(
        n4066) );
  OAI22_X1 U2894 ( .A1(n19844), .A2(n19771), .B1(n20633), .B2(n20503), .ZN(
        n4067) );
  OAI22_X1 U2895 ( .A1(n19844), .A2(n19772), .B1(n20636), .B2(n20504), .ZN(
        n4068) );
  OAI22_X1 U2896 ( .A1(n19844), .A2(n19773), .B1(n20639), .B2(n20504), .ZN(
        n4069) );
  OAI22_X1 U2897 ( .A1(n19844), .A2(n19774), .B1(n20642), .B2(n20503), .ZN(
        n4070) );
  OAI22_X1 U2898 ( .A1(n19844), .A2(n19775), .B1(n20645), .B2(n20500), .ZN(
        n4071) );
  OAI22_X1 U2899 ( .A1(n19844), .A2(n19776), .B1(n20648), .B2(n20499), .ZN(
        n4072) );
  OAI22_X1 U2900 ( .A1(n19844), .A2(n19777), .B1(n20651), .B2(n20502), .ZN(
        n4073) );
  OAI22_X1 U2901 ( .A1(n19844), .A2(n19778), .B1(n20654), .B2(n20501), .ZN(
        n4074) );
  OAI22_X1 U2902 ( .A1(n5126), .A2(n19848), .B1(n20562), .B2(n20516), .ZN(
        n4107) );
  OAI22_X1 U2903 ( .A1(n5127), .A2(n19848), .B1(n20565), .B2(n20515), .ZN(
        n4108) );
  OAI22_X1 U2904 ( .A1(n5128), .A2(n19848), .B1(n20568), .B2(n20516), .ZN(
        n4109) );
  OAI22_X1 U2905 ( .A1(n5129), .A2(n19848), .B1(n20571), .B2(n20518), .ZN(
        n4110) );
  OAI22_X1 U2906 ( .A1(n5130), .A2(n19848), .B1(n20574), .B2(n20516), .ZN(
        n4111) );
  OAI22_X1 U2907 ( .A1(n5131), .A2(n19848), .B1(n20577), .B2(n20521), .ZN(
        n4112) );
  OAI22_X1 U2908 ( .A1(n5132), .A2(n19848), .B1(n20580), .B2(n20517), .ZN(
        n4113) );
  OAI22_X1 U2909 ( .A1(n5133), .A2(n19848), .B1(n20583), .B2(n20518), .ZN(
        n4114) );
  OAI22_X1 U2910 ( .A1(n5134), .A2(n19848), .B1(n20586), .B2(n20518), .ZN(
        n4115) );
  OAI22_X1 U2911 ( .A1(n5135), .A2(n19848), .B1(n20589), .B2(n20520), .ZN(
        n4116) );
  OAI22_X1 U2912 ( .A1(n5136), .A2(n19848), .B1(n20592), .B2(n20519), .ZN(
        n4117) );
  OAI22_X1 U2913 ( .A1(n5137), .A2(n19848), .B1(n20595), .B2(n20520), .ZN(
        n4118) );
  OAI22_X1 U2914 ( .A1(n5138), .A2(n19849), .B1(n20598), .B2(n20517), .ZN(
        n4119) );
  OAI22_X1 U2915 ( .A1(n5139), .A2(n19849), .B1(n20601), .B2(n20518), .ZN(
        n4120) );
  OAI22_X1 U2916 ( .A1(n5140), .A2(n19849), .B1(n20604), .B2(n20517), .ZN(
        n4121) );
  OAI22_X1 U2917 ( .A1(n5141), .A2(n19849), .B1(n20607), .B2(n20519), .ZN(
        n4122) );
  OAI22_X1 U2918 ( .A1(n5142), .A2(n19849), .B1(n20610), .B2(n20519), .ZN(
        n4123) );
  OAI22_X1 U2919 ( .A1(n5143), .A2(n19849), .B1(n20613), .B2(n20520), .ZN(
        n4124) );
  OAI22_X1 U2920 ( .A1(n5144), .A2(n19849), .B1(n20616), .B2(n20520), .ZN(
        n4125) );
  OAI22_X1 U2921 ( .A1(n5145), .A2(n19849), .B1(n20619), .B2(n20516), .ZN(
        n4126) );
  OAI22_X1 U2922 ( .A1(n5146), .A2(n19849), .B1(n20622), .B2(n20519), .ZN(
        n4127) );
  OAI22_X1 U2923 ( .A1(n5147), .A2(n19849), .B1(n20625), .B2(n20522), .ZN(
        n4128) );
  OAI22_X1 U2924 ( .A1(n5148), .A2(n19849), .B1(n20628), .B2(n20522), .ZN(
        n4129) );
  OAI22_X1 U2925 ( .A1(n5149), .A2(n19849), .B1(n20631), .B2(n20521), .ZN(
        n4130) );
  OAI22_X1 U2926 ( .A1(n5150), .A2(n19850), .B1(n20634), .B2(n20521), .ZN(
        n4131) );
  OAI22_X1 U2927 ( .A1(n4889), .A2(n19850), .B1(n20637), .B2(n20522), .ZN(
        n4132) );
  OAI22_X1 U2928 ( .A1(n4890), .A2(n19850), .B1(n20640), .B2(n20522), .ZN(
        n4133) );
  OAI22_X1 U2929 ( .A1(n4891), .A2(n19850), .B1(n20643), .B2(n20521), .ZN(
        n4134) );
  OAI22_X1 U2930 ( .A1(n4892), .A2(n19850), .B1(n20646), .B2(n20515), .ZN(
        n4135) );
  OAI22_X1 U2931 ( .A1(n4893), .A2(n19850), .B1(n20649), .B2(n20515), .ZN(
        n4136) );
  OAI22_X1 U2932 ( .A1(n4894), .A2(n19850), .B1(n20652), .B2(n20515), .ZN(
        n4137) );
  OAI22_X1 U2933 ( .A1(n4895), .A2(n19850), .B1(n20655), .B2(n20517), .ZN(
        n4138) );
  OAI22_X1 U2934 ( .A1(n8657), .A2(n19863), .B1(n20561), .B2(n19893), .ZN(
        n4267) );
  OAI22_X1 U2935 ( .A1(n8658), .A2(n19863), .B1(n20564), .B2(n19894), .ZN(
        n4268) );
  OAI22_X1 U2936 ( .A1(n8659), .A2(n19863), .B1(n20567), .B2(n19894), .ZN(
        n4269) );
  OAI22_X1 U2937 ( .A1(n8660), .A2(n19863), .B1(n20570), .B2(n19895), .ZN(
        n4270) );
  OAI22_X1 U2938 ( .A1(n8661), .A2(n19863), .B1(n20573), .B2(n19893), .ZN(
        n4271) );
  OAI22_X1 U2939 ( .A1(n8662), .A2(n19863), .B1(n20576), .B2(n19895), .ZN(
        n4272) );
  OAI22_X1 U2940 ( .A1(n8663), .A2(n19863), .B1(n20579), .B2(n19894), .ZN(
        n4273) );
  OAI22_X1 U2941 ( .A1(n8664), .A2(n19863), .B1(n20582), .B2(n19895), .ZN(
        n4274) );
  OAI22_X1 U2942 ( .A1(n8671), .A2(n19863), .B1(n20585), .B2(n19893), .ZN(
        n4275) );
  OAI22_X1 U2943 ( .A1(n8665), .A2(n19863), .B1(n20588), .B2(n19893), .ZN(
        n4276) );
  OAI22_X1 U2944 ( .A1(n8666), .A2(n19863), .B1(n20591), .B2(n19894), .ZN(
        n4277) );
  OAI22_X1 U2945 ( .A1(n8672), .A2(n19863), .B1(n20594), .B2(n19894), .ZN(
        n4278) );
  OAI22_X1 U2946 ( .A1(n8673), .A2(n19864), .B1(n20597), .B2(n19895), .ZN(
        n4279) );
  OAI22_X1 U2947 ( .A1(n8674), .A2(n19864), .B1(n20600), .B2(n19893), .ZN(
        n4280) );
  OAI22_X1 U2948 ( .A1(n8675), .A2(n19864), .B1(n20603), .B2(n19895), .ZN(
        n4281) );
  OAI22_X1 U2949 ( .A1(n8667), .A2(n19864), .B1(n20606), .B2(n19894), .ZN(
        n4282) );
  OAI22_X1 U2950 ( .A1(n8668), .A2(n19864), .B1(n20609), .B2(n19895), .ZN(
        n4283) );
  OAI22_X1 U2951 ( .A1(n8676), .A2(n19864), .B1(n20612), .B2(n19893), .ZN(
        n4284) );
  OAI22_X1 U2952 ( .A1(n8669), .A2(n19864), .B1(n20615), .B2(n19893), .ZN(
        n4285) );
  OAI22_X1 U2953 ( .A1(n8670), .A2(n19864), .B1(n20618), .B2(n19894), .ZN(
        n4286) );
  OAI22_X1 U2954 ( .A1(n8677), .A2(n19864), .B1(n20621), .B2(n19894), .ZN(
        n4287) );
  OAI22_X1 U2955 ( .A1(n8678), .A2(n19864), .B1(n20624), .B2(n19895), .ZN(
        n4288) );
  OAI22_X1 U2956 ( .A1(n8679), .A2(n19864), .B1(n20627), .B2(n19893), .ZN(
        n4289) );
  OAI22_X1 U2957 ( .A1(n8680), .A2(n19864), .B1(n20630), .B2(n19895), .ZN(
        n4290) );
  OAI22_X1 U2958 ( .A1(n8681), .A2(n19865), .B1(n20633), .B2(n19894), .ZN(
        n4291) );
  OAI22_X1 U2959 ( .A1(n8682), .A2(n19865), .B1(n20636), .B2(n19895), .ZN(
        n4292) );
  OAI22_X1 U2960 ( .A1(n8686), .A2(n19865), .B1(n20639), .B2(n19893), .ZN(
        n4293) );
  OAI22_X1 U2961 ( .A1(n8683), .A2(n19865), .B1(n20642), .B2(n19893), .ZN(
        n4294) );
  OAI22_X1 U2962 ( .A1(n8684), .A2(n19865), .B1(n20645), .B2(n19894), .ZN(
        n4295) );
  OAI22_X1 U2963 ( .A1(n8687), .A2(n19865), .B1(n20648), .B2(n19894), .ZN(
        n4296) );
  OAI22_X1 U2964 ( .A1(n8688), .A2(n19865), .B1(n20651), .B2(n19895), .ZN(
        n4297) );
  OAI22_X1 U2965 ( .A1(n8685), .A2(n19865), .B1(n20654), .B2(n19893), .ZN(
        n4298) );
  OAI22_X1 U2966 ( .A1(n4843), .A2(n20551), .B1(n20561), .B2(n20559), .ZN(
        n4331) );
  OAI22_X1 U2967 ( .A1(n4844), .A2(n20550), .B1(n20564), .B2(n20559), .ZN(
        n4332) );
  OAI22_X1 U2968 ( .A1(n4845), .A2(n20551), .B1(n20567), .B2(n20559), .ZN(
        n4333) );
  OAI22_X1 U2969 ( .A1(n4846), .A2(n20550), .B1(n20570), .B2(n20559), .ZN(
        n4334) );
  OAI22_X1 U2970 ( .A1(n4847), .A2(n20551), .B1(n20573), .B2(n20558), .ZN(
        n4335) );
  OAI22_X1 U2971 ( .A1(n4848), .A2(n20550), .B1(n20576), .B2(n20558), .ZN(
        n4336) );
  OAI22_X1 U2972 ( .A1(n4849), .A2(n20551), .B1(n20579), .B2(n20558), .ZN(
        n4337) );
  OAI22_X1 U2973 ( .A1(n4850), .A2(n20550), .B1(n20582), .B2(n20558), .ZN(
        n4338) );
  OAI22_X1 U2974 ( .A1(n4851), .A2(n20551), .B1(n20585), .B2(n20557), .ZN(
        n4339) );
  OAI22_X1 U2975 ( .A1(n4852), .A2(n20551), .B1(n20588), .B2(n20557), .ZN(
        n4340) );
  OAI22_X1 U2976 ( .A1(n4853), .A2(n20551), .B1(n20591), .B2(n20557), .ZN(
        n4341) );
  OAI22_X1 U2977 ( .A1(n4854), .A2(n20551), .B1(n20594), .B2(n20557), .ZN(
        n4342) );
  OAI22_X1 U2978 ( .A1(n4855), .A2(n20551), .B1(n20597), .B2(n20556), .ZN(
        n4343) );
  OAI22_X1 U2979 ( .A1(n4856), .A2(n20551), .B1(n20600), .B2(n20556), .ZN(
        n4344) );
  OAI22_X1 U2980 ( .A1(n4857), .A2(n20551), .B1(n20603), .B2(n20556), .ZN(
        n4345) );
  OAI22_X1 U2981 ( .A1(n4858), .A2(n20551), .B1(n20606), .B2(n20556), .ZN(
        n4346) );
  OAI22_X1 U2982 ( .A1(n4859), .A2(n20551), .B1(n20609), .B2(n20555), .ZN(
        n4347) );
  OAI22_X1 U2983 ( .A1(n4860), .A2(n20551), .B1(n20612), .B2(n20555), .ZN(
        n4348) );
  OAI22_X1 U2984 ( .A1(n4861), .A2(n20551), .B1(n20615), .B2(n20555), .ZN(
        n4349) );
  OAI22_X1 U2985 ( .A1(n4862), .A2(n20551), .B1(n20618), .B2(n20555), .ZN(
        n4350) );
  OAI22_X1 U2986 ( .A1(n4863), .A2(n20550), .B1(n20621), .B2(n20554), .ZN(
        n4351) );
  OAI22_X1 U2987 ( .A1(n4864), .A2(n20550), .B1(n20624), .B2(n20554), .ZN(
        n4352) );
  OAI22_X1 U2988 ( .A1(n4865), .A2(n20550), .B1(n20627), .B2(n20554), .ZN(
        n4353) );
  OAI22_X1 U2989 ( .A1(n4866), .A2(n20550), .B1(n20630), .B2(n20554), .ZN(
        n4354) );
  OAI22_X1 U2990 ( .A1(n4867), .A2(n20550), .B1(n20633), .B2(n20553), .ZN(
        n4355) );
  OAI22_X1 U2991 ( .A1(n4868), .A2(n20550), .B1(n20636), .B2(n20553), .ZN(
        n4356) );
  OAI22_X1 U2992 ( .A1(n4869), .A2(n20550), .B1(n20639), .B2(n20553), .ZN(
        n4357) );
  OAI22_X1 U2993 ( .A1(n4870), .A2(n20550), .B1(n20642), .B2(n20553), .ZN(
        n4358) );
  OAI22_X1 U2994 ( .A1(n4871), .A2(n20550), .B1(n20645), .B2(n20552), .ZN(
        n4359) );
  OAI22_X1 U2995 ( .A1(n4872), .A2(n20550), .B1(n20648), .B2(n20552), .ZN(
        n4360) );
  OAI22_X1 U2996 ( .A1(n4873), .A2(n20550), .B1(n20651), .B2(n20552), .ZN(
        n4361) );
  OAI22_X1 U2997 ( .A1(n4874), .A2(n20550), .B1(n20654), .B2(n20552), .ZN(
        n4362) );
  AND3_X1 U2998 ( .A1(ADD_WR[0]), .A2(n1260), .A3(n1586), .ZN(n1447) );
  AND3_X1 U2999 ( .A1(ADD_WR[3]), .A2(ADD_WR[0]), .A3(n1586), .ZN(n1658) );
  AND3_X1 U3000 ( .A1(ADD_WR[3]), .A2(ADD_WR[0]), .A3(n1149), .ZN(n1298) );
  AND3_X1 U3001 ( .A1(n1440), .A2(n1441), .A3(ENABLE), .ZN(n1149) );
  AND3_X1 U3002 ( .A1(n1440), .A2(ADD_WR[4]), .A3(ENABLE), .ZN(n1586) );
  OAI21_X1 U3003 ( .B1(n4396), .B2(n20678), .A(ENABLE), .ZN(n4397) );
  OAI21_X1 U3004 ( .B1(n4398), .B2(n20678), .A(ENABLE), .ZN(n4399) );
  OAI21_X1 U3005 ( .B1(n4400), .B2(n20678), .A(ENABLE), .ZN(n4401) );
  OAI21_X1 U3006 ( .B1(n4402), .B2(n20678), .A(ENABLE), .ZN(n4403) );
  OAI21_X1 U3007 ( .B1(n4404), .B2(n20677), .A(ENABLE), .ZN(n4405) );
  OAI21_X1 U3008 ( .B1(n4406), .B2(n20677), .A(ENABLE), .ZN(n4407) );
  OAI21_X1 U3009 ( .B1(n4408), .B2(n20677), .A(ENABLE), .ZN(n4409) );
  OAI21_X1 U3010 ( .B1(n4410), .B2(n20677), .A(ENABLE), .ZN(n4411) );
  OAI21_X1 U3011 ( .B1(n4412), .B2(n20676), .A(ENABLE), .ZN(n4413) );
  OAI21_X1 U3012 ( .B1(n4414), .B2(n20676), .A(ENABLE), .ZN(n4415) );
  OAI21_X1 U3013 ( .B1(n4416), .B2(n20676), .A(ENABLE), .ZN(n4417) );
  OAI21_X1 U3014 ( .B1(n4418), .B2(n20676), .A(ENABLE), .ZN(n4419) );
  OAI21_X1 U3015 ( .B1(n4420), .B2(n20675), .A(ENABLE), .ZN(n4421) );
  OAI21_X1 U3016 ( .B1(n4422), .B2(n20675), .A(ENABLE), .ZN(n4423) );
  OAI21_X1 U3017 ( .B1(n4424), .B2(n20675), .A(ENABLE), .ZN(n4425) );
  OAI21_X1 U3018 ( .B1(n4426), .B2(n20675), .A(ENABLE), .ZN(n4427) );
  OAI21_X1 U3019 ( .B1(n4428), .B2(n20674), .A(ENABLE), .ZN(n4429) );
  OAI21_X1 U3020 ( .B1(n4430), .B2(n20674), .A(ENABLE), .ZN(n4431) );
  OAI21_X1 U3021 ( .B1(n4432), .B2(n20674), .A(ENABLE), .ZN(n4433) );
  OAI21_X1 U3022 ( .B1(n4434), .B2(n20674), .A(ENABLE), .ZN(n4435) );
  OAI21_X1 U3023 ( .B1(n4436), .B2(n20673), .A(ENABLE), .ZN(n4437) );
  OAI21_X1 U3024 ( .B1(n4438), .B2(n20673), .A(ENABLE), .ZN(n4439) );
  OAI21_X1 U3025 ( .B1(n4440), .B2(n20673), .A(ENABLE), .ZN(n4441) );
  OAI21_X1 U3026 ( .B1(n4442), .B2(n20673), .A(ENABLE), .ZN(n4443) );
  OAI21_X1 U3027 ( .B1(n4444), .B2(n20672), .A(ENABLE), .ZN(n4445) );
  OAI21_X1 U3028 ( .B1(n4446), .B2(n20672), .A(ENABLE), .ZN(n4447) );
  OAI21_X1 U3029 ( .B1(n4448), .B2(n20672), .A(ENABLE), .ZN(n4449) );
  OAI21_X1 U3030 ( .B1(n4450), .B2(n20672), .A(ENABLE), .ZN(n4451) );
  OAI21_X1 U3031 ( .B1(n4452), .B2(n20671), .A(ENABLE), .ZN(n4453) );
  OAI21_X1 U3032 ( .B1(n4454), .B2(n20671), .A(ENABLE), .ZN(n4455) );
  OAI21_X1 U3033 ( .B1(n4456), .B2(n20671), .A(ENABLE), .ZN(n4457) );
  OAI21_X1 U3034 ( .B1(n4458), .B2(n20671), .A(ENABLE), .ZN(n4459) );
  OAI22_X1 U3035 ( .A1(n4972), .A2(n20130), .B1(n18907), .B2(n20137), .ZN(
        n2167) );
  OAI22_X1 U3036 ( .A1(n4973), .A2(n20130), .B1(n18908), .B2(n20136), .ZN(
        n2142) );
  OAI22_X1 U3037 ( .A1(n4974), .A2(n20130), .B1(n18909), .B2(n20138), .ZN(
        n2117) );
  OAI22_X1 U3038 ( .A1(n4975), .A2(n20125), .B1(n18910), .B2(n20136), .ZN(
        n2092) );
  OAI22_X1 U3039 ( .A1(n4977), .A2(n20128), .B1(n18911), .B2(n20133), .ZN(
        n2067) );
  OAI22_X1 U3040 ( .A1(n4882), .A2(n20126), .B1(n18912), .B2(n20138), .ZN(
        n2042) );
  OAI22_X1 U3041 ( .A1(n4883), .A2(n20129), .B1(n18913), .B2(n20138), .ZN(
        n2017) );
  OAI22_X1 U3042 ( .A1(n4884), .A2(n20130), .B1(n18914), .B2(n20138), .ZN(
        n1992) );
  AND3_X1 U3043 ( .A1(ADD_WR[3]), .A2(n1437), .A3(n1586), .ZN(n1655) );
  INV_X1 U3044 ( .A(RD1), .ZN(n5722) );
  OAI21_X1 U3045 ( .B1(n3083), .B2(n19884), .A(ENABLE), .ZN(n3084) );
  OAI21_X1 U3046 ( .B1(n3089), .B2(n19885), .A(ENABLE), .ZN(n3090) );
  OAI21_X1 U3047 ( .B1(n3095), .B2(n19884), .A(ENABLE), .ZN(n3096) );
  OAI21_X1 U3048 ( .B1(n3101), .B2(n19885), .A(ENABLE), .ZN(n3102) );
  OAI21_X1 U3049 ( .B1(n3107), .B2(n19886), .A(ENABLE), .ZN(n3108) );
  OAI21_X1 U3050 ( .B1(n3113), .B2(n19884), .A(ENABLE), .ZN(n3114) );
  OAI21_X1 U3051 ( .B1(n3119), .B2(n19886), .A(ENABLE), .ZN(n3120) );
  OAI21_X1 U3052 ( .B1(n3149), .B2(n19885), .A(ENABLE), .ZN(n3150) );
  OAI21_X1 U3053 ( .B1(n3167), .B2(n19884), .A(ENABLE), .ZN(n3168) );
  OAI21_X1 U3054 ( .B1(n3173), .B2(n19885), .A(ENABLE), .ZN(n3174) );
  OAI21_X1 U3055 ( .B1(n3179), .B2(n19886), .A(ENABLE), .ZN(n3180) );
  OAI21_X1 U3056 ( .B1(n3185), .B2(n19886), .A(ENABLE), .ZN(n3186) );
  OAI21_X1 U3057 ( .B1(n3191), .B2(n19884), .A(ENABLE), .ZN(n3192) );
  OAI21_X1 U3058 ( .B1(n3197), .B2(n19885), .A(ENABLE), .ZN(n3198) );
  OAI21_X1 U3059 ( .B1(n3227), .B2(n19886), .A(ENABLE), .ZN(n3228) );
  OAI21_X1 U3060 ( .B1(n3239), .B2(n19884), .A(ENABLE), .ZN(n3240) );
  OAI21_X1 U3061 ( .B1(n3245), .B2(n19885), .A(ENABLE), .ZN(n3246) );
  OAI21_X1 U3062 ( .B1(n3251), .B2(n19886), .A(ENABLE), .ZN(n3252) );
  OAI21_X1 U3063 ( .B1(n3125), .B2(n19887), .A(ENABLE), .ZN(n3126) );
  OAI21_X1 U3064 ( .B1(n3131), .B2(n19887), .A(ENABLE), .ZN(n3132) );
  OAI21_X1 U3065 ( .B1(n3137), .B2(n19888), .A(ENABLE), .ZN(n3138) );
  OAI21_X1 U3066 ( .B1(n3155), .B2(n19888), .A(ENABLE), .ZN(n3156) );
  OAI21_X1 U3067 ( .B1(n3203), .B2(n19887), .A(ENABLE), .ZN(n3204) );
  OAI21_X1 U3068 ( .B1(n3209), .B2(n19888), .A(ENABLE), .ZN(n3210) );
  OAI21_X1 U3069 ( .B1(n3221), .B2(n19887), .A(ENABLE), .ZN(n3222) );
  OAI21_X1 U3070 ( .B1(n3233), .B2(n19887), .A(ENABLE), .ZN(n3234) );
  OAI21_X1 U3071 ( .B1(n3257), .B2(n19888), .A(ENABLE), .ZN(n3258) );
  OAI21_X1 U3072 ( .B1(n3263), .B2(n19888), .A(ENABLE), .ZN(n3264) );
  OAI21_X1 U3073 ( .B1(n3143), .B2(n19889), .A(ENABLE), .ZN(n3144) );
  OAI21_X1 U3074 ( .B1(n3161), .B2(n19889), .A(ENABLE), .ZN(n3162) );
  OAI21_X1 U3075 ( .B1(n3215), .B2(n19889), .A(ENABLE), .ZN(n3216) );
  OAI21_X1 U3076 ( .B1(n3269), .B2(n19889), .A(ENABLE), .ZN(n3270) );
  INV_X1 U3077 ( .A(RD2), .ZN(n2646) );
  NOR2_X1 U3078 ( .A1(ADD_WR[3]), .A2(ADD_WR[0]), .ZN(n1150) );
  INV_X1 U3079 ( .A(ADD_WR[1]), .ZN(n1727) );
  INV_X1 U3080 ( .A(ADD_WR[2]), .ZN(n1796) );
  INV_X1 U3081 ( .A(ADD_WR[0]), .ZN(n1437) );
  INV_X1 U3082 ( .A(ADD_WR[3]), .ZN(n1260) );
  INV_X1 U3083 ( .A(ADD_WR[4]), .ZN(n1441) );
  INV_X1 U3084 ( .A(RESET), .ZN(n20758) );
  NAND3_X1 U3085 ( .A1(n2646), .A2(n20746), .A3(ENABLE), .ZN(n19866) );
  NAND3_X1 U3086 ( .A1(n2646), .A2(n20746), .A3(ENABLE), .ZN(n19867) );
  NAND3_X1 U3087 ( .A1(n5722), .A2(n20746), .A3(ENABLE), .ZN(n19874) );
  NAND3_X1 U3088 ( .A1(n5722), .A2(n20746), .A3(ENABLE), .ZN(n19875) );
  NAND3_X1 U3089 ( .A1(n5684), .A2(n5722), .A3(ENABLE), .ZN(n19882) );
  NAND3_X1 U3090 ( .A1(n5684), .A2(n5722), .A3(ENABLE), .ZN(n19883) );
  INV_X1 U3091 ( .A(n2745), .ZN(n19896) );
  INV_X1 U3092 ( .A(n19896), .ZN(n19897) );
  INV_X1 U3093 ( .A(n19896), .ZN(n19898) );
  INV_X1 U3094 ( .A(n19896), .ZN(n19899) );
  INV_X1 U3095 ( .A(n19896), .ZN(n19900) );
  INV_X1 U3096 ( .A(n19896), .ZN(n19901) );
  INV_X1 U3097 ( .A(n19896), .ZN(n19902) );
  INV_X1 U3098 ( .A(n19896), .ZN(n19903) );
  INV_X1 U3099 ( .A(n2746), .ZN(n19904) );
  INV_X1 U3100 ( .A(n19904), .ZN(n19905) );
  INV_X1 U3101 ( .A(n19904), .ZN(n19906) );
  INV_X1 U3102 ( .A(n19904), .ZN(n19907) );
  INV_X1 U3103 ( .A(n19904), .ZN(n19908) );
  INV_X1 U3104 ( .A(n19904), .ZN(n19909) );
  INV_X1 U3105 ( .A(n19904), .ZN(n19910) );
  INV_X1 U3106 ( .A(n19904), .ZN(n19911) );
  INV_X1 U3107 ( .A(n19912), .ZN(n19914) );
  INV_X1 U3108 ( .A(n19912), .ZN(n19915) );
  INV_X1 U3109 ( .A(n19912), .ZN(n19916) );
  INV_X1 U3110 ( .A(n19913), .ZN(n19917) );
  INV_X1 U3111 ( .A(n19913), .ZN(n19918) );
  INV_X1 U3112 ( .A(n19913), .ZN(n19919) );
  INV_X1 U3113 ( .A(n19920), .ZN(n19922) );
  INV_X1 U3114 ( .A(n19920), .ZN(n19923) );
  INV_X1 U3115 ( .A(n19920), .ZN(n19924) );
  INV_X1 U3116 ( .A(n19921), .ZN(n19925) );
  INV_X1 U3117 ( .A(n19921), .ZN(n19926) );
  INV_X1 U3118 ( .A(n19921), .ZN(n19927) );
  INV_X1 U3119 ( .A(n2740), .ZN(n19928) );
  INV_X1 U3120 ( .A(n19928), .ZN(n19929) );
  INV_X1 U3121 ( .A(n19928), .ZN(n19930) );
  INV_X1 U3122 ( .A(n19928), .ZN(n19931) );
  INV_X1 U3123 ( .A(n19928), .ZN(n19932) );
  INV_X1 U3124 ( .A(n19928), .ZN(n19933) );
  INV_X1 U3125 ( .A(n19928), .ZN(n19934) );
  INV_X1 U3126 ( .A(n19928), .ZN(n19935) );
  INV_X1 U3127 ( .A(n2741), .ZN(n19936) );
  INV_X1 U3128 ( .A(n19936), .ZN(n19937) );
  INV_X1 U3129 ( .A(n19936), .ZN(n19938) );
  INV_X1 U3130 ( .A(n19936), .ZN(n19939) );
  INV_X1 U3131 ( .A(n19936), .ZN(n19940) );
  INV_X1 U3132 ( .A(n19936), .ZN(n19941) );
  INV_X1 U3133 ( .A(n19936), .ZN(n19942) );
  INV_X1 U3134 ( .A(n19936), .ZN(n19943) );
  INV_X1 U3135 ( .A(n19944), .ZN(n19946) );
  INV_X1 U3136 ( .A(n19944), .ZN(n19947) );
  INV_X1 U3137 ( .A(n19944), .ZN(n19948) );
  INV_X1 U3138 ( .A(n19945), .ZN(n19949) );
  INV_X1 U3139 ( .A(n19945), .ZN(n19950) );
  INV_X1 U3140 ( .A(n19945), .ZN(n19951) );
  INV_X1 U3141 ( .A(n19952), .ZN(n19953) );
  INV_X1 U3142 ( .A(n19952), .ZN(n19954) );
  INV_X1 U3143 ( .A(n19952), .ZN(n19955) );
  INV_X1 U3144 ( .A(n19952), .ZN(n19956) );
  INV_X1 U3145 ( .A(n19952), .ZN(n19957) );
  INV_X1 U3146 ( .A(n19952), .ZN(n19958) );
  INV_X1 U3147 ( .A(n19952), .ZN(n19959) );
  INV_X1 U3148 ( .A(n2729), .ZN(n19960) );
  INV_X1 U3149 ( .A(n19960), .ZN(n19961) );
  INV_X1 U3150 ( .A(n19960), .ZN(n19962) );
  INV_X1 U3151 ( .A(n19960), .ZN(n19963) );
  INV_X1 U3152 ( .A(n19960), .ZN(n19964) );
  INV_X1 U3153 ( .A(n19960), .ZN(n19965) );
  INV_X1 U3154 ( .A(n19960), .ZN(n19966) );
  INV_X1 U3155 ( .A(n19960), .ZN(n19967) );
  INV_X1 U3156 ( .A(n19968), .ZN(n19969) );
  INV_X1 U3157 ( .A(n19968), .ZN(n19970) );
  INV_X1 U3158 ( .A(n19968), .ZN(n19971) );
  INV_X1 U3159 ( .A(n19968), .ZN(n19972) );
  INV_X1 U3160 ( .A(n19968), .ZN(n19973) );
  INV_X1 U3161 ( .A(n19968), .ZN(n19974) );
  INV_X1 U3162 ( .A(n19968), .ZN(n19975) );
  INV_X1 U3163 ( .A(n19976), .ZN(n19977) );
  INV_X1 U3164 ( .A(n19976), .ZN(n19978) );
  INV_X1 U3165 ( .A(n19976), .ZN(n19979) );
  INV_X1 U3166 ( .A(n19976), .ZN(n19980) );
  INV_X1 U3167 ( .A(n19976), .ZN(n19981) );
  INV_X1 U3168 ( .A(n19976), .ZN(n19982) );
  INV_X1 U3169 ( .A(n19976), .ZN(n19983) );
  INV_X1 U3170 ( .A(n2737), .ZN(n19984) );
  INV_X1 U3171 ( .A(n19984), .ZN(n19985) );
  INV_X1 U3172 ( .A(n19984), .ZN(n19986) );
  INV_X1 U3173 ( .A(n19984), .ZN(n19987) );
  INV_X1 U3174 ( .A(n19984), .ZN(n19988) );
  INV_X1 U3175 ( .A(n19984), .ZN(n19989) );
  INV_X1 U3176 ( .A(n19984), .ZN(n19990) );
  INV_X1 U3177 ( .A(n19984), .ZN(n19991) );
  INV_X1 U3178 ( .A(n2738), .ZN(n19992) );
  INV_X1 U3179 ( .A(n19992), .ZN(n19993) );
  INV_X1 U3180 ( .A(n19992), .ZN(n19994) );
  INV_X1 U3181 ( .A(n19992), .ZN(n19995) );
  INV_X1 U3182 ( .A(n19992), .ZN(n19996) );
  INV_X1 U3183 ( .A(n19992), .ZN(n19997) );
  INV_X1 U3184 ( .A(n19992), .ZN(n19998) );
  INV_X1 U3185 ( .A(n19992), .ZN(n19999) );
  INV_X1 U3186 ( .A(n20000), .ZN(n20001) );
  INV_X1 U3187 ( .A(n20000), .ZN(n20002) );
  INV_X1 U3188 ( .A(n20000), .ZN(n20003) );
  INV_X1 U3189 ( .A(n20000), .ZN(n20004) );
  INV_X1 U3190 ( .A(n20000), .ZN(n20005) );
  INV_X1 U3191 ( .A(n20000), .ZN(n20006) );
  INV_X1 U3192 ( .A(n20000), .ZN(n20007) );
  INV_X1 U3193 ( .A(n20008), .ZN(n20009) );
  INV_X1 U3194 ( .A(n20008), .ZN(n20010) );
  INV_X1 U3195 ( .A(n20008), .ZN(n20011) );
  INV_X1 U3196 ( .A(n20008), .ZN(n20012) );
  INV_X1 U3197 ( .A(n20008), .ZN(n20013) );
  INV_X1 U3198 ( .A(n20008), .ZN(n20014) );
  INV_X1 U3199 ( .A(n20008), .ZN(n20015) );
  INV_X1 U3200 ( .A(n20016), .ZN(n20017) );
  INV_X1 U3201 ( .A(n20016), .ZN(n20018) );
  INV_X1 U3202 ( .A(n20016), .ZN(n20019) );
  INV_X1 U3203 ( .A(n20016), .ZN(n20020) );
  INV_X1 U3204 ( .A(n20016), .ZN(n20021) );
  INV_X1 U3205 ( .A(n20016), .ZN(n20022) );
  INV_X1 U3206 ( .A(n20016), .ZN(n20023) );
  INV_X1 U3207 ( .A(n20024), .ZN(n20025) );
  INV_X1 U3208 ( .A(n20024), .ZN(n20026) );
  INV_X1 U3209 ( .A(n20024), .ZN(n20027) );
  INV_X1 U3210 ( .A(n20024), .ZN(n20028) );
  INV_X1 U3211 ( .A(n20024), .ZN(n20029) );
  INV_X1 U3212 ( .A(n20024), .ZN(n20030) );
  INV_X1 U3213 ( .A(n20024), .ZN(n20031) );
  INV_X1 U3214 ( .A(n2726), .ZN(n20032) );
  INV_X1 U3215 ( .A(n20032), .ZN(n20033) );
  INV_X1 U3216 ( .A(n20032), .ZN(n20034) );
  INV_X1 U3217 ( .A(n20032), .ZN(n20035) );
  INV_X1 U3218 ( .A(n20032), .ZN(n20036) );
  INV_X1 U3219 ( .A(n20032), .ZN(n20037) );
  INV_X1 U3220 ( .A(n20032), .ZN(n20038) );
  INV_X1 U3221 ( .A(n20032), .ZN(n20039) );
  INV_X1 U3222 ( .A(n20049), .ZN(n20050) );
  INV_X1 U3223 ( .A(n20049), .ZN(n20051) );
  INV_X1 U3224 ( .A(n20049), .ZN(n20052) );
  INV_X1 U3225 ( .A(n20049), .ZN(n20053) );
  INV_X1 U3226 ( .A(n20049), .ZN(n20054) );
  INV_X1 U3227 ( .A(n20049), .ZN(n20055) );
  INV_X1 U3228 ( .A(n20049), .ZN(n20056) );
  INV_X1 U3229 ( .A(n2720), .ZN(n20057) );
  INV_X1 U3230 ( .A(n20057), .ZN(n20058) );
  INV_X1 U3231 ( .A(n20057), .ZN(n20059) );
  INV_X1 U3232 ( .A(n20057), .ZN(n20060) );
  INV_X1 U3233 ( .A(n20057), .ZN(n20061) );
  INV_X1 U3234 ( .A(n20057), .ZN(n20062) );
  INV_X1 U3235 ( .A(n20057), .ZN(n20063) );
  INV_X1 U3236 ( .A(n20057), .ZN(n20064) );
  INV_X1 U3237 ( .A(n2721), .ZN(n20065) );
  INV_X1 U3238 ( .A(n20065), .ZN(n20066) );
  INV_X1 U3239 ( .A(n20065), .ZN(n20067) );
  INV_X1 U3240 ( .A(n20065), .ZN(n20068) );
  INV_X1 U3241 ( .A(n20065), .ZN(n20069) );
  INV_X1 U3242 ( .A(n20065), .ZN(n20070) );
  INV_X1 U3243 ( .A(n20065), .ZN(n20071) );
  INV_X1 U3244 ( .A(n20065), .ZN(n20072) );
  INV_X1 U3245 ( .A(n20074), .ZN(n20075) );
  INV_X1 U3246 ( .A(n20073), .ZN(n20076) );
  INV_X1 U3247 ( .A(n20073), .ZN(n20077) );
  INV_X1 U3248 ( .A(n20073), .ZN(n20078) );
  INV_X1 U3249 ( .A(n20074), .ZN(n20079) );
  INV_X1 U3250 ( .A(n20074), .ZN(n20080) );
  INV_X1 U3251 ( .A(n1887), .ZN(n20107) );
  INV_X1 U3252 ( .A(n1887), .ZN(n20108) );
  INV_X1 U3253 ( .A(n20108), .ZN(n20109) );
  INV_X1 U3254 ( .A(n20108), .ZN(n20110) );
  INV_X1 U3255 ( .A(n20107), .ZN(n20111) );
  INV_X1 U3256 ( .A(n20107), .ZN(n20112) );
  INV_X1 U3257 ( .A(n20108), .ZN(n20113) );
  INV_X1 U3258 ( .A(n20108), .ZN(n20114) );
  INV_X1 U3259 ( .A(n1889), .ZN(n20115) );
  INV_X1 U3260 ( .A(n20115), .ZN(n20116) );
  INV_X1 U3261 ( .A(n20115), .ZN(n20117) );
  INV_X1 U3262 ( .A(n20115), .ZN(n20118) );
  INV_X1 U3263 ( .A(n20115), .ZN(n20119) );
  INV_X1 U3264 ( .A(n20115), .ZN(n20120) );
  INV_X1 U3265 ( .A(n20115), .ZN(n20121) );
  INV_X1 U3266 ( .A(n20115), .ZN(n20122) );
  INV_X1 U3267 ( .A(n20123), .ZN(n20124) );
  INV_X1 U3268 ( .A(n20123), .ZN(n20125) );
  INV_X1 U3269 ( .A(n20123), .ZN(n20126) );
  INV_X1 U3270 ( .A(n20123), .ZN(n20127) );
  INV_X1 U3271 ( .A(n20123), .ZN(n20128) );
  INV_X1 U3272 ( .A(n20123), .ZN(n20129) );
  INV_X1 U3273 ( .A(n20123), .ZN(n20130) );
  INV_X1 U3274 ( .A(n20131), .ZN(n20132) );
  INV_X1 U3275 ( .A(n20131), .ZN(n20133) );
  INV_X1 U3276 ( .A(n20131), .ZN(n20134) );
  INV_X1 U3277 ( .A(n20131), .ZN(n20135) );
  INV_X1 U3278 ( .A(n20131), .ZN(n20136) );
  INV_X1 U3279 ( .A(n20131), .ZN(n20137) );
  INV_X1 U3280 ( .A(n20131), .ZN(n20138) );
  INV_X1 U3281 ( .A(n1882), .ZN(n20139) );
  INV_X1 U3282 ( .A(n20139), .ZN(n20140) );
  INV_X1 U3283 ( .A(n20139), .ZN(n20141) );
  INV_X1 U3284 ( .A(n20139), .ZN(n20142) );
  INV_X1 U3285 ( .A(n20139), .ZN(n20143) );
  INV_X1 U3286 ( .A(n20139), .ZN(n20144) );
  INV_X1 U3287 ( .A(n20139), .ZN(n20145) );
  INV_X1 U3288 ( .A(n20139), .ZN(n20146) );
  INV_X1 U3289 ( .A(n1883), .ZN(n20147) );
  INV_X1 U3290 ( .A(n1883), .ZN(n20148) );
  INV_X1 U3291 ( .A(n20147), .ZN(n20149) );
  INV_X1 U3292 ( .A(n20147), .ZN(n20150) );
  INV_X1 U3293 ( .A(n20147), .ZN(n20151) );
  INV_X1 U3294 ( .A(n20148), .ZN(n20152) );
  INV_X1 U3295 ( .A(n20148), .ZN(n20153) );
  INV_X1 U3296 ( .A(n20148), .ZN(n20154) );
  INV_X1 U3297 ( .A(n20155), .ZN(n20156) );
  INV_X1 U3298 ( .A(n20155), .ZN(n20157) );
  INV_X1 U3299 ( .A(n20155), .ZN(n20158) );
  INV_X1 U3300 ( .A(n20155), .ZN(n20159) );
  INV_X1 U3301 ( .A(n20155), .ZN(n20160) );
  INV_X1 U3302 ( .A(n20155), .ZN(n20161) );
  INV_X1 U3303 ( .A(n20155), .ZN(n20162) );
  INV_X1 U3304 ( .A(n20163), .ZN(n20164) );
  INV_X1 U3305 ( .A(n20163), .ZN(n20165) );
  INV_X1 U3306 ( .A(n20163), .ZN(n20166) );
  INV_X1 U3307 ( .A(n20163), .ZN(n20167) );
  INV_X1 U3308 ( .A(n20163), .ZN(n20168) );
  INV_X1 U3309 ( .A(n20163), .ZN(n20169) );
  INV_X1 U3310 ( .A(n20163), .ZN(n20170) );
  INV_X1 U3311 ( .A(n1871), .ZN(n20171) );
  INV_X1 U3312 ( .A(n20171), .ZN(n20172) );
  INV_X1 U3313 ( .A(n20171), .ZN(n20173) );
  INV_X1 U3314 ( .A(n20171), .ZN(n20174) );
  INV_X1 U3315 ( .A(n20171), .ZN(n20175) );
  INV_X1 U3316 ( .A(n20171), .ZN(n20176) );
  INV_X1 U3317 ( .A(n20171), .ZN(n20177) );
  INV_X1 U3318 ( .A(n20171), .ZN(n20178) );
  INV_X1 U3319 ( .A(n20179), .ZN(n20180) );
  INV_X1 U3320 ( .A(n20179), .ZN(n20181) );
  INV_X1 U3321 ( .A(n20179), .ZN(n20182) );
  INV_X1 U3322 ( .A(n20179), .ZN(n20183) );
  INV_X1 U3323 ( .A(n20179), .ZN(n20184) );
  INV_X1 U3324 ( .A(n20179), .ZN(n20185) );
  INV_X1 U3325 ( .A(n20179), .ZN(n20186) );
  INV_X1 U3326 ( .A(n20187), .ZN(n20188) );
  INV_X1 U3327 ( .A(n20187), .ZN(n20189) );
  INV_X1 U3328 ( .A(n20187), .ZN(n20190) );
  INV_X1 U3329 ( .A(n20187), .ZN(n20191) );
  INV_X1 U3330 ( .A(n20187), .ZN(n20192) );
  INV_X1 U3331 ( .A(n20187), .ZN(n20193) );
  INV_X1 U3332 ( .A(n20187), .ZN(n20194) );
  INV_X1 U3333 ( .A(n1880), .ZN(n20195) );
  INV_X1 U3334 ( .A(n20195), .ZN(n20196) );
  INV_X1 U3335 ( .A(n20195), .ZN(n20197) );
  INV_X1 U3336 ( .A(n20195), .ZN(n20198) );
  INV_X1 U3337 ( .A(n20195), .ZN(n20199) );
  INV_X1 U3338 ( .A(n20195), .ZN(n20200) );
  INV_X1 U3339 ( .A(n20195), .ZN(n20201) );
  INV_X1 U3340 ( .A(n20195), .ZN(n20202) );
  INV_X1 U3341 ( .A(n1881), .ZN(n20203) );
  INV_X1 U3342 ( .A(n1881), .ZN(n20204) );
  INV_X1 U3343 ( .A(n20203), .ZN(n20205) );
  INV_X1 U3344 ( .A(n20204), .ZN(n20206) );
  INV_X1 U3345 ( .A(n20203), .ZN(n20207) );
  INV_X1 U3346 ( .A(n20203), .ZN(n20208) );
  INV_X1 U3347 ( .A(n20204), .ZN(n20209) );
  INV_X1 U3348 ( .A(n20204), .ZN(n20210) );
  INV_X1 U3349 ( .A(n20211), .ZN(n20212) );
  INV_X1 U3350 ( .A(n20211), .ZN(n20213) );
  INV_X1 U3351 ( .A(n20211), .ZN(n20214) );
  INV_X1 U3352 ( .A(n20211), .ZN(n20215) );
  INV_X1 U3353 ( .A(n20211), .ZN(n20216) );
  INV_X1 U3354 ( .A(n20211), .ZN(n20217) );
  INV_X1 U3355 ( .A(n20211), .ZN(n20218) );
  INV_X1 U3356 ( .A(n20220), .ZN(n20221) );
  INV_X1 U3357 ( .A(n20219), .ZN(n20222) );
  INV_X1 U3358 ( .A(n20219), .ZN(n20223) );
  INV_X1 U3359 ( .A(n20219), .ZN(n20224) );
  INV_X1 U3360 ( .A(n20220), .ZN(n20225) );
  INV_X1 U3361 ( .A(n20220), .ZN(n20226) );
  INV_X1 U3362 ( .A(n20227), .ZN(n20228) );
  INV_X1 U3363 ( .A(n20227), .ZN(n20229) );
  INV_X1 U3364 ( .A(n20227), .ZN(n20230) );
  INV_X1 U3365 ( .A(n20227), .ZN(n20231) );
  INV_X1 U3366 ( .A(n20227), .ZN(n20232) );
  INV_X1 U3367 ( .A(n20227), .ZN(n20233) );
  INV_X1 U3368 ( .A(n20227), .ZN(n20234) );
  INV_X1 U3369 ( .A(n20235), .ZN(n20236) );
  INV_X1 U3370 ( .A(n20235), .ZN(n20237) );
  INV_X1 U3371 ( .A(n20235), .ZN(n20238) );
  INV_X1 U3372 ( .A(n20235), .ZN(n20239) );
  INV_X1 U3373 ( .A(n20235), .ZN(n20240) );
  INV_X1 U3374 ( .A(n20235), .ZN(n20241) );
  INV_X1 U3375 ( .A(n20235), .ZN(n20242) );
  INV_X1 U3376 ( .A(n1868), .ZN(n20243) );
  INV_X1 U3377 ( .A(n20243), .ZN(n20244) );
  INV_X1 U3378 ( .A(n20243), .ZN(n20245) );
  INV_X1 U3379 ( .A(n20243), .ZN(n20246) );
  INV_X1 U3380 ( .A(n20243), .ZN(n20247) );
  INV_X1 U3381 ( .A(n20243), .ZN(n20248) );
  INV_X1 U3382 ( .A(n20243), .ZN(n20249) );
  INV_X1 U3383 ( .A(n20243), .ZN(n20250) );
  INV_X1 U3384 ( .A(n1870), .ZN(n20251) );
  INV_X1 U3385 ( .A(n20251), .ZN(n20252) );
  INV_X1 U3386 ( .A(n20251), .ZN(n20253) );
  INV_X1 U3387 ( .A(n20251), .ZN(n20254) );
  INV_X1 U3388 ( .A(n20251), .ZN(n20255) );
  INV_X1 U3389 ( .A(n20251), .ZN(n20256) );
  INV_X1 U3390 ( .A(n20251), .ZN(n20257) );
  INV_X1 U3391 ( .A(n20251), .ZN(n20258) );
  INV_X1 U3392 ( .A(n20259), .ZN(n20260) );
  INV_X1 U3393 ( .A(n20259), .ZN(n20261) );
  INV_X1 U3394 ( .A(n20259), .ZN(n20262) );
  INV_X1 U3395 ( .A(n20259), .ZN(n20263) );
  INV_X1 U3396 ( .A(n20259), .ZN(n20264) );
  INV_X1 U3397 ( .A(n20259), .ZN(n20265) );
  INV_X1 U3398 ( .A(n20259), .ZN(n20266) );
  INV_X1 U3399 ( .A(n1863), .ZN(n20269) );
  INV_X1 U3400 ( .A(n20269), .ZN(n20270) );
  INV_X1 U3401 ( .A(n20269), .ZN(n20271) );
  INV_X1 U3402 ( .A(n20269), .ZN(n20272) );
  INV_X1 U3403 ( .A(n20269), .ZN(n20273) );
  INV_X1 U3404 ( .A(n20269), .ZN(n20274) );
  INV_X1 U3405 ( .A(n20269), .ZN(n20275) );
  INV_X1 U3406 ( .A(n20269), .ZN(n20276) );
  INV_X1 U3407 ( .A(n1864), .ZN(n20277) );
  INV_X1 U3408 ( .A(n1864), .ZN(n20278) );
  INV_X1 U3409 ( .A(n20277), .ZN(n20279) );
  INV_X1 U3410 ( .A(n20278), .ZN(n20280) );
  INV_X1 U3411 ( .A(n20277), .ZN(n20281) );
  INV_X1 U3412 ( .A(n20278), .ZN(n20282) );
  INV_X1 U3413 ( .A(n20278), .ZN(n20283) );
  INV_X1 U3414 ( .A(n20277), .ZN(n20284) );
  INV_X1 U3415 ( .A(n20298), .ZN(n20299) );
  INV_X1 U3416 ( .A(n20298), .ZN(n20300) );
  INV_X1 U3417 ( .A(n20298), .ZN(n20301) );
  INV_X1 U3418 ( .A(n20298), .ZN(n20302) );
  INV_X1 U3419 ( .A(n20298), .ZN(n20303) );
  INV_X1 U3420 ( .A(n20298), .ZN(n20304) );
  INV_X1 U3421 ( .A(n20298), .ZN(n20305) );
  INV_X1 U3422 ( .A(n20321), .ZN(n20322) );
  INV_X1 U3423 ( .A(n20320), .ZN(n20323) );
  INV_X1 U3424 ( .A(n20320), .ZN(n20324) );
  INV_X1 U3425 ( .A(n20321), .ZN(n20325) );
  INV_X1 U3426 ( .A(n20321), .ZN(n20326) );
  INV_X1 U3427 ( .A(n20321), .ZN(n20327) );
  INV_X1 U3428 ( .A(n20321), .ZN(n20328) );
  INV_X1 U3429 ( .A(n20330), .ZN(n20331) );
  INV_X1 U3430 ( .A(n20329), .ZN(n20332) );
  INV_X1 U3431 ( .A(n20329), .ZN(n20333) );
  INV_X1 U3432 ( .A(n20330), .ZN(n20334) );
  INV_X1 U3433 ( .A(n20330), .ZN(n20335) );
  INV_X1 U3434 ( .A(n20330), .ZN(n20336) );
  INV_X1 U3435 ( .A(n20330), .ZN(n20337) );
  INV_X1 U3436 ( .A(n20338), .ZN(n20340) );
  INV_X1 U3437 ( .A(n20338), .ZN(n20341) );
  INV_X1 U3438 ( .A(n20338), .ZN(n20342) );
  INV_X1 U3439 ( .A(n20338), .ZN(n20343) );
  INV_X1 U3440 ( .A(n20338), .ZN(n20344) );
  INV_X1 U3441 ( .A(n20338), .ZN(n20345) );
  INV_X1 U3442 ( .A(n20339), .ZN(n20346) );
  INV_X1 U3443 ( .A(n20348), .ZN(n20349) );
  INV_X1 U3444 ( .A(n20347), .ZN(n20350) );
  INV_X1 U3445 ( .A(n20347), .ZN(n20351) );
  INV_X1 U3446 ( .A(n20348), .ZN(n20352) );
  INV_X1 U3447 ( .A(n20348), .ZN(n20353) );
  INV_X1 U3448 ( .A(n20348), .ZN(n20354) );
  INV_X1 U3449 ( .A(n20348), .ZN(n20355) );
  INV_X1 U3450 ( .A(n20356), .ZN(n20358) );
  INV_X1 U3451 ( .A(n20356), .ZN(n20359) );
  INV_X1 U3452 ( .A(n20356), .ZN(n20360) );
  INV_X1 U3453 ( .A(n20356), .ZN(n20361) );
  INV_X1 U3454 ( .A(n20356), .ZN(n20362) );
  INV_X1 U3455 ( .A(n20356), .ZN(n20363) );
  INV_X1 U3456 ( .A(n20357), .ZN(n20364) );
  INV_X1 U3457 ( .A(n20366), .ZN(n20367) );
  INV_X1 U3458 ( .A(n20365), .ZN(n20368) );
  INV_X1 U3459 ( .A(n20365), .ZN(n20369) );
  INV_X1 U3460 ( .A(n20366), .ZN(n20370) );
  INV_X1 U3461 ( .A(n20366), .ZN(n20371) );
  INV_X1 U3462 ( .A(n20366), .ZN(n20372) );
  INV_X1 U3463 ( .A(n20366), .ZN(n20373) );
  INV_X1 U3464 ( .A(n20374), .ZN(n20375) );
  INV_X1 U3465 ( .A(n20374), .ZN(n20376) );
  INV_X1 U3466 ( .A(n20374), .ZN(n20377) );
  INV_X1 U3467 ( .A(n20374), .ZN(n20378) );
  INV_X1 U3468 ( .A(n20374), .ZN(n20379) );
  INV_X1 U3469 ( .A(n20374), .ZN(n20380) );
  INV_X1 U3470 ( .A(n20374), .ZN(n20381) );
  INV_X1 U3471 ( .A(n20374), .ZN(n20382) );
  INV_X1 U3472 ( .A(n20384), .ZN(n20385) );
  INV_X1 U3473 ( .A(n20383), .ZN(n20386) );
  INV_X1 U3474 ( .A(n20383), .ZN(n20387) );
  INV_X1 U3475 ( .A(n20384), .ZN(n20388) );
  INV_X1 U3476 ( .A(n20384), .ZN(n20389) );
  INV_X1 U3477 ( .A(n20384), .ZN(n20390) );
  INV_X1 U3478 ( .A(n20384), .ZN(n20391) );
  INV_X1 U3479 ( .A(n20393), .ZN(n20394) );
  INV_X1 U3480 ( .A(n20392), .ZN(n20395) );
  INV_X1 U3481 ( .A(n20392), .ZN(n20396) );
  INV_X1 U3482 ( .A(n20393), .ZN(n20397) );
  INV_X1 U3483 ( .A(n20393), .ZN(n20398) );
  INV_X1 U3484 ( .A(n20393), .ZN(n20399) );
  INV_X1 U3485 ( .A(n20393), .ZN(n20400) );
  INV_X1 U3486 ( .A(n20401), .ZN(n20403) );
  INV_X1 U3487 ( .A(n20401), .ZN(n20404) );
  INV_X1 U3488 ( .A(n20401), .ZN(n20405) );
  INV_X1 U3489 ( .A(n20401), .ZN(n20406) );
  INV_X1 U3490 ( .A(n20401), .ZN(n20407) );
  INV_X1 U3491 ( .A(n20401), .ZN(n20408) );
  INV_X1 U3492 ( .A(n20402), .ZN(n20409) );
  INV_X1 U3493 ( .A(n20411), .ZN(n20412) );
  INV_X1 U3494 ( .A(n20410), .ZN(n20413) );
  INV_X1 U3495 ( .A(n20410), .ZN(n20414) );
  INV_X1 U3496 ( .A(n20411), .ZN(n20415) );
  INV_X1 U3497 ( .A(n20411), .ZN(n20416) );
  INV_X1 U3498 ( .A(n20411), .ZN(n20417) );
  INV_X1 U3499 ( .A(n20411), .ZN(n20418) );
  INV_X1 U3500 ( .A(n20419), .ZN(n20420) );
  INV_X1 U3501 ( .A(n20419), .ZN(n20421) );
  INV_X1 U3502 ( .A(n20419), .ZN(n20422) );
  INV_X1 U3503 ( .A(n20419), .ZN(n20423) );
  INV_X1 U3504 ( .A(n20419), .ZN(n20424) );
  INV_X1 U3505 ( .A(n20419), .ZN(n20425) );
  INV_X1 U3506 ( .A(n20419), .ZN(n20426) );
  INV_X1 U3507 ( .A(n20419), .ZN(n20427) );
  INV_X1 U3508 ( .A(n20429), .ZN(n20430) );
  INV_X1 U3509 ( .A(n20428), .ZN(n20431) );
  INV_X1 U3510 ( .A(n20428), .ZN(n20432) );
  INV_X1 U3511 ( .A(n20429), .ZN(n20433) );
  INV_X1 U3512 ( .A(n20429), .ZN(n20434) );
  INV_X1 U3513 ( .A(n20429), .ZN(n20435) );
  INV_X1 U3514 ( .A(n20429), .ZN(n20436) );
  INV_X1 U3515 ( .A(n20438), .ZN(n20439) );
  INV_X1 U3516 ( .A(n20437), .ZN(n20440) );
  INV_X1 U3517 ( .A(n20437), .ZN(n20441) );
  INV_X1 U3518 ( .A(n20438), .ZN(n20442) );
  INV_X1 U3519 ( .A(n20438), .ZN(n20443) );
  INV_X1 U3520 ( .A(n20438), .ZN(n20444) );
  INV_X1 U3521 ( .A(n20438), .ZN(n20445) );
  INV_X1 U3522 ( .A(n20446), .ZN(n20447) );
  INV_X1 U3523 ( .A(n20446), .ZN(n20448) );
  INV_X1 U3524 ( .A(n20446), .ZN(n20449) );
  INV_X1 U3525 ( .A(n20446), .ZN(n20450) );
  INV_X1 U3526 ( .A(n20446), .ZN(n20451) );
  INV_X1 U3527 ( .A(n20446), .ZN(n20452) );
  INV_X1 U3528 ( .A(n20446), .ZN(n20453) );
  INV_X1 U3529 ( .A(n20446), .ZN(n20454) );
  INV_X1 U3530 ( .A(n20455), .ZN(n20456) );
  INV_X1 U3531 ( .A(n20455), .ZN(n20457) );
  INV_X1 U3532 ( .A(n20455), .ZN(n20458) );
  INV_X1 U3533 ( .A(n20455), .ZN(n20459) );
  INV_X1 U3534 ( .A(n20455), .ZN(n20460) );
  INV_X1 U3535 ( .A(n20455), .ZN(n20461) );
  INV_X1 U3536 ( .A(n20455), .ZN(n20462) );
  INV_X1 U3537 ( .A(n20455), .ZN(n20463) );
  INV_X1 U3538 ( .A(n20464), .ZN(n20465) );
  INV_X1 U3539 ( .A(n20464), .ZN(n20466) );
  INV_X1 U3540 ( .A(n20464), .ZN(n20467) );
  INV_X1 U3541 ( .A(n20464), .ZN(n20468) );
  INV_X1 U3542 ( .A(n20464), .ZN(n20469) );
  INV_X1 U3543 ( .A(n20464), .ZN(n20470) );
  INV_X1 U3545 ( .A(n20464), .ZN(n20471) );
  INV_X1 U3546 ( .A(n20464), .ZN(n20472) );
  INV_X1 U3547 ( .A(n20481), .ZN(n20482) );
  INV_X1 U3548 ( .A(n20480), .ZN(n20483) );
  INV_X1 U3549 ( .A(n20480), .ZN(n20484) );
  INV_X1 U3550 ( .A(n20481), .ZN(n20485) );
  INV_X1 U3551 ( .A(n20481), .ZN(n20486) );
  INV_X1 U3552 ( .A(n20481), .ZN(n20487) );
  INV_X1 U3553 ( .A(n20481), .ZN(n20488) );
  INV_X1 U3554 ( .A(n20497), .ZN(n20498) );
  INV_X1 U3555 ( .A(n20496), .ZN(n20499) );
  INV_X1 U3556 ( .A(n20496), .ZN(n20500) );
  INV_X1 U3557 ( .A(n20497), .ZN(n20501) );
  INV_X1 U3558 ( .A(n20497), .ZN(n20502) );
  INV_X1 U3559 ( .A(n20497), .ZN(n20503) );
  INV_X1 U3560 ( .A(n20497), .ZN(n20504) );
  INV_X1 U3561 ( .A(n20505), .ZN(n20507) );
  INV_X1 U3562 ( .A(n20505), .ZN(n20508) );
  INV_X1 U3563 ( .A(n20505), .ZN(n20509) );
  INV_X1 U3564 ( .A(n20505), .ZN(n20510) );
  INV_X1 U3565 ( .A(n20505), .ZN(n20511) );
  INV_X1 U3566 ( .A(n20505), .ZN(n20512) );
  INV_X1 U3567 ( .A(n20506), .ZN(n20513) );
  INV_X1 U3568 ( .A(n20514), .ZN(n20515) );
  INV_X1 U3569 ( .A(n20514), .ZN(n20516) );
  INV_X1 U3570 ( .A(n20514), .ZN(n20517) );
  INV_X1 U3571 ( .A(n20514), .ZN(n20518) );
  INV_X1 U3572 ( .A(n20514), .ZN(n20519) );
  INV_X1 U3573 ( .A(n20514), .ZN(n20520) );
  INV_X1 U3574 ( .A(n20514), .ZN(n20521) );
  INV_X1 U3575 ( .A(n20514), .ZN(n20522) );
  INV_X1 U3576 ( .A(n20524), .ZN(n20525) );
  INV_X1 U3577 ( .A(n20523), .ZN(n20526) );
  INV_X1 U3578 ( .A(n20523), .ZN(n20527) );
  INV_X1 U3579 ( .A(n20524), .ZN(n20528) );
  INV_X1 U3580 ( .A(n20524), .ZN(n20529) );
  INV_X1 U3581 ( .A(n20524), .ZN(n20530) );
  INV_X1 U3582 ( .A(n20524), .ZN(n20531) );
  CLKBUF_X1 U3583 ( .A(n20756), .Z(n20687) );
  CLKBUF_X1 U3584 ( .A(n20756), .Z(n20688) );
  CLKBUF_X1 U3585 ( .A(n20756), .Z(n20689) );
  CLKBUF_X1 U3586 ( .A(n20756), .Z(n20690) );
  CLKBUF_X1 U3587 ( .A(n20756), .Z(n20691) );
  CLKBUF_X1 U3588 ( .A(n20756), .Z(n20692) );
  CLKBUF_X1 U3589 ( .A(n20755), .Z(n20693) );
  CLKBUF_X1 U3590 ( .A(n20755), .Z(n20694) );
  CLKBUF_X1 U3591 ( .A(n20755), .Z(n20695) );
  CLKBUF_X1 U3592 ( .A(n20755), .Z(n20696) );
  CLKBUF_X1 U3593 ( .A(n20755), .Z(n20697) );
  CLKBUF_X1 U3594 ( .A(n20755), .Z(n20698) );
  CLKBUF_X1 U3595 ( .A(n20754), .Z(n20699) );
  CLKBUF_X1 U3596 ( .A(n20754), .Z(n20700) );
  CLKBUF_X1 U3597 ( .A(n20754), .Z(n20701) );
  CLKBUF_X1 U3598 ( .A(n20754), .Z(n20702) );
  CLKBUF_X1 U3599 ( .A(n20754), .Z(n20703) );
  CLKBUF_X1 U3600 ( .A(n20754), .Z(n20704) );
  CLKBUF_X1 U3601 ( .A(n20753), .Z(n20705) );
  CLKBUF_X1 U3602 ( .A(n20753), .Z(n20706) );
  CLKBUF_X1 U3603 ( .A(n20753), .Z(n20707) );
  CLKBUF_X1 U3604 ( .A(n20753), .Z(n20708) );
  CLKBUF_X1 U3605 ( .A(n20753), .Z(n20709) );
  CLKBUF_X1 U3606 ( .A(n20753), .Z(n20710) );
  CLKBUF_X1 U3607 ( .A(n20752), .Z(n20711) );
  CLKBUF_X1 U3608 ( .A(n20752), .Z(n20712) );
  CLKBUF_X1 U3609 ( .A(n20752), .Z(n20713) );
  CLKBUF_X1 U3610 ( .A(n20752), .Z(n20714) );
  CLKBUF_X1 U3611 ( .A(n20752), .Z(n20715) );
  CLKBUF_X1 U3612 ( .A(n20752), .Z(n20716) );
  CLKBUF_X1 U3613 ( .A(n20751), .Z(n20717) );
  CLKBUF_X1 U3614 ( .A(n20751), .Z(n20718) );
  CLKBUF_X1 U3615 ( .A(n20751), .Z(n20719) );
  CLKBUF_X1 U3616 ( .A(n20751), .Z(n20720) );
  CLKBUF_X1 U3617 ( .A(n20751), .Z(n20721) );
  CLKBUF_X1 U3635 ( .A(n20751), .Z(n20722) );
  CLKBUF_X1 U3636 ( .A(n20750), .Z(n20723) );
  CLKBUF_X1 U3637 ( .A(n20750), .Z(n20724) );
  CLKBUF_X1 U3638 ( .A(n20750), .Z(n20725) );
  CLKBUF_X1 U3639 ( .A(n20750), .Z(n20726) );
  CLKBUF_X1 U3640 ( .A(n20750), .Z(n20727) );
  CLKBUF_X1 U3641 ( .A(n20750), .Z(n20728) );
  CLKBUF_X1 U3642 ( .A(n20749), .Z(n20729) );
  CLKBUF_X1 U3643 ( .A(n20749), .Z(n20730) );
  CLKBUF_X1 U3644 ( .A(n20749), .Z(n20731) );
  CLKBUF_X1 U3645 ( .A(n20749), .Z(n20732) );
  CLKBUF_X1 U3646 ( .A(n20749), .Z(n20733) );
  CLKBUF_X1 U3647 ( .A(n20749), .Z(n20734) );
  CLKBUF_X1 U3648 ( .A(n20748), .Z(n20735) );
  CLKBUF_X1 U3649 ( .A(n20748), .Z(n20736) );
  CLKBUF_X1 U3650 ( .A(n20748), .Z(n20737) );
  CLKBUF_X1 U3651 ( .A(n20748), .Z(n20738) );
  CLKBUF_X1 U3652 ( .A(n20748), .Z(n20739) );
  CLKBUF_X1 U3653 ( .A(n20748), .Z(n20740) );
  CLKBUF_X1 U3654 ( .A(n20747), .Z(n20741) );
  CLKBUF_X1 U3655 ( .A(n20747), .Z(n20742) );
  CLKBUF_X1 U3656 ( .A(n20747), .Z(n20743) );
  CLKBUF_X1 U3657 ( .A(n20747), .Z(n20744) );
  CLKBUF_X1 U3658 ( .A(n20747), .Z(n20745) );
  CLKBUF_X1 U3659 ( .A(n20747), .Z(n20746) );
endmodule


module mux41N_Nbit5 ( in3, in2, in1, in0, sel, Y );
  input [4:0] in3;
  input [4:0] in2;
  input [4:0] in1;
  input [4:0] in0;
  input [1:0] sel;
  output [4:0] Y;
  wire   \outmux[2][4] , \outmux[2][3] , \outmux[2][2] , \outmux[2][1] ,
         \outmux[2][0] , \outmux[1][4] , \outmux[1][3] , \outmux[1][2] ,
         \outmux[1][1] , \outmux[1][0] ;
  tri   [1:0] sel;

  mux21N_N5_35 row1_1 ( .in1(in1), .in0(in0), .S(sel[0]), .U({\outmux[1][4] , 
        \outmux[1][3] , \outmux[1][2] , \outmux[1][1] , \outmux[1][0] }) );
  mux21N_N5_34 row1_2 ( .in1(in3), .in0(in2), .S(sel[0]), .U({\outmux[2][4] , 
        \outmux[2][3] , \outmux[2][2] , \outmux[2][1] , \outmux[2][0] }) );
  mux21N_N5_33 row2_1 ( .in1({\outmux[2][4] , \outmux[2][3] , \outmux[2][2] , 
        \outmux[2][1] , \outmux[2][0] }), .in0({\outmux[1][4] , \outmux[1][3] , 
        \outmux[1][2] , \outmux[1][1] , \outmux[1][0] }), .S(sel[1]), .U(Y) );
endmodule


module mux21N_N5_36 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;

  tri   S;

  MUX21_571 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_570 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_569 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_568 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_567 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module mux21N_N5_8 ( in1, in0, S, U );
  input [4:0] in1;
  input [4:0] in0;
  output [4:0] U;
  input S;

  tri   S;

  MUX21_576 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(S), .Y(U[0]) );
  MUX21_575 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(S), .Y(U[1]) );
  MUX21_574 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(S), .Y(U[2]) );
  MUX21_573 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(S), .Y(U[3]) );
  MUX21_572 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(S), .Y(U[4]) );
endmodule


module FD_EN_437 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module RegEn_Nbit32_10 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;
  wire   n21, n22, n23, n24;
  assign n21 = Reset;

  FD_EN_335 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[0]) );
  FD_EN_334 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[1]) );
  FD_EN_333 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[2]) );
  FD_EN_332 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[3]) );
  FD_EN_331 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[4]) );
  FD_EN_330 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[5]) );
  FD_EN_329 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[6]) );
  FD_EN_328 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[7]) );
  FD_EN_327 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[8]) );
  FD_EN_326 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[9]) );
  FD_EN_325 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[10]) );
  FD_EN_324 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[11]) );
  FD_EN_323 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[12]) );
  FD_EN_322 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[13]) );
  FD_EN_321 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[14]) );
  FD_EN_320 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[15]) );
  FD_EN_319 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[16]) );
  FD_EN_318 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[17]) );
  FD_EN_317 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[18]) );
  FD_EN_316 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[19]) );
  FD_EN_315 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[20]) );
  FD_EN_314 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[21]) );
  FD_EN_313 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[22]) );
  FD_EN_312 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[23]) );
  FD_EN_311 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[24]) );
  FD_EN_310 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[25]) );
  FD_EN_309 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[26]) );
  FD_EN_308 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[27]) );
  FD_EN_307 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[28]) );
  FD_EN_306 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[29]) );
  FD_EN_305 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[30]) );
  FD_EN_304 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[31]) );
  BUF_X1 U1 ( .A(n21), .Z(n22) );
  BUF_X1 U2 ( .A(n21), .Z(n23) );
  BUF_X1 U3 ( .A(n21), .Z(n24) );
endmodule


module RegEn_Nbit32_11 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;
  wire   n21, n22, n23, n24;
  assign n21 = Reset;

  FD_EN_367 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[0]) );
  FD_EN_366 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[1]) );
  FD_EN_365 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[2]) );
  FD_EN_364 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[3]) );
  FD_EN_363 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[4]) );
  FD_EN_362 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[5]) );
  FD_EN_361 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[6]) );
  FD_EN_360 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[7]) );
  FD_EN_359 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[8]) );
  FD_EN_358 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[9]) );
  FD_EN_357 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[10]) );
  FD_EN_356 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(n22), .EN(EN), .Q(U[11]) );
  FD_EN_355 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[12]) );
  FD_EN_354 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[13]) );
  FD_EN_353 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[14]) );
  FD_EN_352 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[15]) );
  FD_EN_351 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[16]) );
  FD_EN_350 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[17]) );
  FD_EN_349 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[18]) );
  FD_EN_348 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[19]) );
  FD_EN_347 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[20]) );
  FD_EN_346 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[21]) );
  FD_EN_345 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[22]) );
  FD_EN_344 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(n23), .EN(EN), .Q(U[23]) );
  FD_EN_343 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[24]) );
  FD_EN_342 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[25]) );
  FD_EN_341 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[26]) );
  FD_EN_340 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[27]) );
  FD_EN_339 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[28]) );
  FD_EN_338 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[29]) );
  FD_EN_337 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[30]) );
  FD_EN_336 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(n24), .EN(EN), .Q(U[31]) );
  BUF_X1 U1 ( .A(n21), .Z(n22) );
  BUF_X1 U2 ( .A(n21), .Z(n23) );
  BUF_X1 U3 ( .A(n21), .Z(n24) );
endmodule


module RegEn_Nbit32_12 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;


  FD_EN_399 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_398 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_397 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_396 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_395 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
  FD_EN_394 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[5]) );
  FD_EN_393 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[6]) );
  FD_EN_392 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[7]) );
  FD_EN_391 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[8]) );
  FD_EN_390 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[9]) );
  FD_EN_389 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[10])
         );
  FD_EN_388 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[11])
         );
  FD_EN_387 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[12])
         );
  FD_EN_386 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[13])
         );
  FD_EN_385 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[14])
         );
  FD_EN_384 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[15])
         );
  FD_EN_383 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[16])
         );
  FD_EN_382 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[17])
         );
  FD_EN_381 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[18])
         );
  FD_EN_380 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[19])
         );
  FD_EN_379 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[20])
         );
  FD_EN_378 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[21])
         );
  FD_EN_377 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[22])
         );
  FD_EN_376 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[23])
         );
  FD_EN_375 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[24])
         );
  FD_EN_374 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[25])
         );
  FD_EN_373 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[26])
         );
  FD_EN_372 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[27])
         );
  FD_EN_371 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[28])
         );
  FD_EN_370 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[29])
         );
  FD_EN_369 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[30])
         );
  FD_EN_368 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[31])
         );
endmodule


module FD_EN_438 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n4, n2, n3;

  DFF_X1 Q_reg ( .D(n4), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n2), .ZN(n4) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module mux21N_N30_1 ( in1, in0, S, U );
  input [29:0] in1;
  input [29:0] in0;
  output [29:0] U;
  input S;
  wire   n21, n22, n23, n24;
  assign n21 = S;

  MUX21_606 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n22), .Y(U[0]) );
  MUX21_605 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n22), .Y(U[1]) );
  MUX21_604 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n22), .Y(U[2]) );
  MUX21_603 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n22), .Y(U[3]) );
  MUX21_602 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n22), .Y(U[4]) );
  MUX21_601 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n22), .Y(U[5]) );
  MUX21_600 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n22), .Y(U[6]) );
  MUX21_599 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n22), .Y(U[7]) );
  MUX21_598 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n22), .Y(U[8]) );
  MUX21_597 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n22), .Y(U[9]) );
  MUX21_596 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n22), .Y(U[10]) );
  MUX21_595 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n22), .Y(U[11]) );
  MUX21_594 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n23), .Y(U[12]) );
  MUX21_593 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n23), .Y(U[13]) );
  MUX21_592 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n23), .Y(U[14]) );
  MUX21_591 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n23), .Y(U[15]) );
  MUX21_590 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n23), .Y(U[16]) );
  MUX21_589 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n23), .Y(U[17]) );
  MUX21_588 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n23), .Y(U[18]) );
  MUX21_587 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n23), .Y(U[19]) );
  MUX21_586 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n23), .Y(U[20]) );
  MUX21_585 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n23), .Y(U[21]) );
  MUX21_584 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n23), .Y(U[22]) );
  MUX21_583 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n23), .Y(U[23]) );
  MUX21_582 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n24), .Y(U[24]) );
  MUX21_581 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n24), .Y(U[25]) );
  MUX21_580 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n24), .Y(U[26]) );
  MUX21_579 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n24), .Y(U[27]) );
  MUX21_578 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n24), .Y(U[28]) );
  MUX21_577 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n24), .Y(U[29]) );
  BUF_X1 U1 ( .A(n21), .Z(n22) );
  BUF_X1 U2 ( .A(n21), .Z(n23) );
  BUF_X1 U3 ( .A(n21), .Z(n24) );
endmodule


module mux21N_N30_0 ( in1, in0, S, U );
  input [29:0] in1;
  input [29:0] in0;
  output [29:0] U;
  input S;
  wire   n24, n25, n26, n27;
  assign n24 = S;

  MUX21_636 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n25), .Y(U[0]) );
  MUX21_635 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n25), .Y(U[1]) );
  MUX21_634 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n25), .Y(U[2]) );
  MUX21_633 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n25), .Y(U[3]) );
  MUX21_632 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n25), .Y(U[4]) );
  MUX21_631 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n25), .Y(U[5]) );
  MUX21_630 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n25), .Y(U[6]) );
  MUX21_629 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n25), .Y(U[7]) );
  MUX21_628 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n25), .Y(U[8]) );
  MUX21_627 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n25), .Y(U[9]) );
  MUX21_626 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n25), .Y(U[10]) );
  MUX21_625 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n25), .Y(U[11]) );
  MUX21_624 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n26), .Y(U[12]) );
  MUX21_623 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n26), .Y(U[13]) );
  MUX21_622 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n26), .Y(U[14]) );
  MUX21_621 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n26), .Y(U[15]) );
  MUX21_620 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n26), .Y(U[16]) );
  MUX21_619 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n26), .Y(U[17]) );
  MUX21_618 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n26), .Y(U[18]) );
  MUX21_617 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n26), .Y(U[19]) );
  MUX21_616 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n26), .Y(U[20]) );
  MUX21_615 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n26), .Y(U[21]) );
  MUX21_614 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n26), .Y(U[22]) );
  MUX21_613 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n26), .Y(U[23]) );
  MUX21_612 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n27), .Y(U[24]) );
  MUX21_611 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n27), .Y(U[25]) );
  MUX21_610 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n27), .Y(U[26]) );
  MUX21_609 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n27), .Y(U[27]) );
  MUX21_608 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n27), .Y(U[28]) );
  MUX21_607 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n27), .Y(U[29]) );
  CLKBUF_X1 U1 ( .A(n24), .Z(n25) );
  CLKBUF_X1 U2 ( .A(n24), .Z(n26) );
  CLKBUF_X1 U3 ( .A(n24), .Z(n27) );
endmodule


module mux21N_N32_13 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   n24, n25, n26, n27;
  assign n24 = S;

  MUX21_668 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n25), .Y(U[0]) );
  MUX21_667 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n25), .Y(U[1]) );
  MUX21_666 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n25), .Y(U[2]) );
  MUX21_665 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n25), .Y(U[3]) );
  MUX21_664 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n25), .Y(U[4]) );
  MUX21_663 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n25), .Y(U[5]) );
  MUX21_662 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n25), .Y(U[6]) );
  MUX21_661 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n25), .Y(U[7]) );
  MUX21_660 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n25), .Y(U[8]) );
  MUX21_659 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n25), .Y(U[9]) );
  MUX21_658 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n25), .Y(U[10]) );
  MUX21_657 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n25), .Y(U[11]) );
  MUX21_656 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n26), .Y(U[12]) );
  MUX21_655 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n26), .Y(U[13]) );
  MUX21_654 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n26), .Y(U[14]) );
  MUX21_653 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n26), .Y(U[15]) );
  MUX21_652 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n26), .Y(U[16]) );
  MUX21_651 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n26), .Y(U[17]) );
  MUX21_650 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n26), .Y(U[18]) );
  MUX21_649 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n26), .Y(U[19]) );
  MUX21_648 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n27), .Y(U[20]) );
  MUX21_647 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n26), .Y(U[21]) );
  MUX21_646 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n26), .Y(U[22]) );
  MUX21_645 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n26), .Y(U[23]) );
  MUX21_644 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n26), .Y(U[24]) );
  MUX21_643 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n27), .Y(U[25]) );
  MUX21_642 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n27), .Y(U[26]) );
  MUX21_641 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n27), .Y(U[27]) );
  MUX21_640 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n27), .Y(U[28]) );
  MUX21_639 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n27), .Y(U[29]) );
  MUX21_638 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n27), .Y(U[30]) );
  MUX21_637 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n27), .Y(U[31]) );
  CLKBUF_X1 U1 ( .A(n24), .Z(n26) );
  CLKBUF_X1 U2 ( .A(n24), .Z(n25) );
  CLKBUF_X1 U3 ( .A(n24), .Z(n27) );
endmodule


module mux21N_N32_14 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   n24, n25, n26, n27;
  assign n24 = S;

  MUX21_700 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n25), .Y(U[0]) );
  MUX21_699 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n25), .Y(U[1]) );
  MUX21_698 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n25), .Y(U[2]) );
  MUX21_697 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n25), .Y(U[3]) );
  MUX21_696 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n25), .Y(U[4]) );
  MUX21_695 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n25), .Y(U[5]) );
  MUX21_694 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n25), .Y(U[6]) );
  MUX21_693 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n25), .Y(U[7]) );
  MUX21_692 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n25), .Y(U[8]) );
  MUX21_691 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n25), .Y(U[9]) );
  MUX21_690 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n25), .Y(U[10]) );
  MUX21_689 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n25), .Y(U[11]) );
  MUX21_688 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n26), .Y(U[12]) );
  MUX21_687 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n26), .Y(U[13]) );
  MUX21_686 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n26), .Y(U[14]) );
  MUX21_685 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n26), .Y(U[15]) );
  MUX21_684 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n26), .Y(U[16]) );
  MUX21_683 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n26), .Y(U[17]) );
  MUX21_682 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n26), .Y(U[18]) );
  MUX21_681 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n26), .Y(U[19]) );
  MUX21_680 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n26), .Y(U[20]) );
  MUX21_679 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n26), .Y(U[21]) );
  MUX21_678 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n26), .Y(U[22]) );
  MUX21_677 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n26), .Y(U[23]) );
  MUX21_676 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n27), .Y(U[24]) );
  MUX21_675 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n27), .Y(U[25]) );
  MUX21_674 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n27), .Y(U[26]) );
  MUX21_673 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n27), .Y(U[27]) );
  MUX21_672 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n27), .Y(U[28]) );
  MUX21_671 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n27), .Y(U[29]) );
  MUX21_670 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n27), .Y(U[30]) );
  MUX21_669 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n27), .Y(U[31]) );
  CLKBUF_X1 U1 ( .A(n24), .Z(n26) );
  CLKBUF_X1 U2 ( .A(n24), .Z(n25) );
  CLKBUF_X1 U3 ( .A(n24), .Z(n27) );
endmodule


module RegEn_Nbit32_0 ( A, Clk, Reset, EN, U );
  input [31:0] A;
  output [31:0] U;
  input Clk, Reset, EN;


  FD_EN_431 FDS_0 ( .D(A[0]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[0]) );
  FD_EN_430 FDS_1 ( .D(A[1]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[1]) );
  FD_EN_429 FDS_2 ( .D(A[2]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[2]) );
  FD_EN_428 FDS_3 ( .D(A[3]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[3]) );
  FD_EN_427 FDS_4 ( .D(A[4]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[4]) );
  FD_EN_426 FDS_5 ( .D(A[5]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[5]) );
  FD_EN_425 FDS_6 ( .D(A[6]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[6]) );
  FD_EN_424 FDS_7 ( .D(A[7]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[7]) );
  FD_EN_423 FDS_8 ( .D(A[8]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[8]) );
  FD_EN_422 FDS_9 ( .D(A[9]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[9]) );
  FD_EN_421 FDS_10 ( .D(A[10]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[10])
         );
  FD_EN_420 FDS_11 ( .D(A[11]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[11])
         );
  FD_EN_419 FDS_12 ( .D(A[12]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[12])
         );
  FD_EN_418 FDS_13 ( .D(A[13]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[13])
         );
  FD_EN_417 FDS_14 ( .D(A[14]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[14])
         );
  FD_EN_416 FDS_15 ( .D(A[15]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[15])
         );
  FD_EN_415 FDS_16 ( .D(A[16]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[16])
         );
  FD_EN_414 FDS_17 ( .D(A[17]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[17])
         );
  FD_EN_413 FDS_18 ( .D(A[18]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[18])
         );
  FD_EN_412 FDS_19 ( .D(A[19]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[19])
         );
  FD_EN_411 FDS_20 ( .D(A[20]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[20])
         );
  FD_EN_410 FDS_21 ( .D(A[21]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[21])
         );
  FD_EN_409 FDS_22 ( .D(A[22]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[22])
         );
  FD_EN_408 FDS_23 ( .D(A[23]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[23])
         );
  FD_EN_407 FDS_24 ( .D(A[24]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[24])
         );
  FD_EN_406 FDS_25 ( .D(A[25]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[25])
         );
  FD_EN_405 FDS_26 ( .D(A[26]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[26])
         );
  FD_EN_404 FDS_27 ( .D(A[27]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[27])
         );
  FD_EN_403 FDS_28 ( .D(A[28]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[28])
         );
  FD_EN_402 FDS_29 ( .D(A[29]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[29])
         );
  FD_EN_401 FDS_30 ( .D(A[30]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[30])
         );
  FD_EN_400 FDS_31 ( .D(A[31]), .Clk(Clk), .RESET(Reset), .EN(EN), .Q(U[31])
         );
endmodule


module MUX21_800 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n4), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n4) );
endmodule


module mux41 ( in3, in2, in1, in0, sel, Y );
  input [1:0] sel;
  input in3, in2, in1, in0;
  output Y;

  wire   [2:1] outmux;
  tri   [1:0] sel;

  MUX21_703 row1_1 ( .in1(in1), .in0(in0), .S(sel[0]), .Y(outmux[1]) );
  MUX21_702 row1_2 ( .in1(in3), .in0(in2), .S(sel[0]), .Y(outmux[2]) );
  MUX21_701 row2_1 ( .in1(outmux[2]), .in0(outmux[1]), .S(sel[1]), .Y(Y) );
endmodule


module FD_EN_0 ( D, Clk, RESET, EN, Q );
  input D, Clk, RESET, EN;
  output Q;
  wire   n5, n2, n3;

  DFF_X1 Q_reg ( .D(n5), .CK(Clk), .Q(Q) );
  NOR2_X1 U3 ( .A1(RESET), .A2(n2), .ZN(n5) );
  AOI22_X1 U4 ( .A1(EN), .A2(D), .B1(n3), .B2(Q), .ZN(n2) );
  INV_X1 U5 ( .A(EN), .ZN(n3) );
endmodule


module AddSubN_Nbit32_0 ( A, B, addnsub, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input addnsub;
  output Cout;

  wire   [31:0] addendB;
  wire   [7:0] Carry;

  SparseTreeCarryGenN_Nbit32_0 STCG ( .A(A), .B(addendB), .Cin(addnsub), 
        .Cout({Cout, Carry}) );
  CarrySumN_Nbit32_0 CSN ( .A(A), .B(addendB), .Ci(Carry), .S(S) );
  XOR2_X1 U1 ( .A(addnsub), .B(B[9]), .Z(addendB[9]) );
  XOR2_X1 U2 ( .A(addnsub), .B(B[8]), .Z(addendB[8]) );
  XOR2_X1 U3 ( .A(addnsub), .B(B[7]), .Z(addendB[7]) );
  XOR2_X1 U4 ( .A(addnsub), .B(B[6]), .Z(addendB[6]) );
  XOR2_X1 U5 ( .A(addnsub), .B(B[5]), .Z(addendB[5]) );
  XOR2_X1 U6 ( .A(addnsub), .B(B[4]), .Z(addendB[4]) );
  XOR2_X1 U7 ( .A(addnsub), .B(B[3]), .Z(addendB[3]) );
  XOR2_X1 U8 ( .A(addnsub), .B(B[31]), .Z(addendB[31]) );
  XOR2_X1 U9 ( .A(addnsub), .B(B[30]), .Z(addendB[30]) );
  XOR2_X1 U10 ( .A(addnsub), .B(B[2]), .Z(addendB[2]) );
  XOR2_X1 U11 ( .A(addnsub), .B(B[29]), .Z(addendB[29]) );
  XOR2_X1 U12 ( .A(addnsub), .B(B[28]), .Z(addendB[28]) );
  XOR2_X1 U13 ( .A(addnsub), .B(B[27]), .Z(addendB[27]) );
  XOR2_X1 U14 ( .A(addnsub), .B(B[26]), .Z(addendB[26]) );
  XOR2_X1 U15 ( .A(addnsub), .B(B[25]), .Z(addendB[25]) );
  XOR2_X1 U16 ( .A(addnsub), .B(B[24]), .Z(addendB[24]) );
  XOR2_X1 U17 ( .A(addnsub), .B(B[23]), .Z(addendB[23]) );
  XOR2_X1 U18 ( .A(addnsub), .B(B[22]), .Z(addendB[22]) );
  XOR2_X1 U19 ( .A(addnsub), .B(B[21]), .Z(addendB[21]) );
  XOR2_X1 U20 ( .A(addnsub), .B(B[20]), .Z(addendB[20]) );
  XOR2_X1 U21 ( .A(addnsub), .B(B[1]), .Z(addendB[1]) );
  XOR2_X1 U22 ( .A(addnsub), .B(B[19]), .Z(addendB[19]) );
  XOR2_X1 U23 ( .A(addnsub), .B(B[18]), .Z(addendB[18]) );
  XOR2_X1 U24 ( .A(addnsub), .B(B[17]), .Z(addendB[17]) );
  XOR2_X1 U25 ( .A(addnsub), .B(B[16]), .Z(addendB[16]) );
  XOR2_X1 U26 ( .A(addnsub), .B(B[15]), .Z(addendB[15]) );
  XOR2_X1 U27 ( .A(addnsub), .B(B[14]), .Z(addendB[14]) );
  XOR2_X1 U28 ( .A(addnsub), .B(B[13]), .Z(addendB[13]) );
  XOR2_X1 U29 ( .A(addnsub), .B(B[12]), .Z(addendB[12]) );
  XOR2_X1 U30 ( .A(addnsub), .B(B[11]), .Z(addendB[11]) );
  XOR2_X1 U31 ( .A(addnsub), .B(B[10]), .Z(addendB[10]) );
  XOR2_X1 U32 ( .A(addnsub), .B(B[0]), .Z(addendB[0]) );
endmodule


module mux21N_N32_15 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   n21, n22, n23, n24;
  assign n21 = S;

  MUX21_735 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n24), .Y(U[0]) );
  MUX21_734 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n22), .Y(U[1]) );
  MUX21_733 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n22), .Y(U[2]) );
  MUX21_732 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n22), .Y(U[3]) );
  MUX21_731 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n22), .Y(U[4]) );
  MUX21_730 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n22), .Y(U[5]) );
  MUX21_729 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n22), .Y(U[6]) );
  MUX21_728 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n22), .Y(U[7]) );
  MUX21_727 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n22), .Y(U[8]) );
  MUX21_726 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n22), .Y(U[9]) );
  MUX21_725 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n22), .Y(U[10]) );
  MUX21_724 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n22), .Y(U[11]) );
  MUX21_723 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n22), .Y(U[12]) );
  MUX21_722 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n23), .Y(U[13]) );
  MUX21_721 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n23), .Y(U[14]) );
  MUX21_720 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n23), .Y(U[15]) );
  MUX21_719 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n23), .Y(U[16]) );
  MUX21_718 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n23), .Y(U[17]) );
  MUX21_717 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n23), .Y(U[18]) );
  MUX21_716 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n23), .Y(U[19]) );
  MUX21_715 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n23), .Y(U[20]) );
  MUX21_714 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n23), .Y(U[21]) );
  MUX21_713 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n23), .Y(U[22]) );
  MUX21_712 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n23), .Y(U[23]) );
  MUX21_711 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n23), .Y(U[24]) );
  MUX21_710 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n24), .Y(U[25]) );
  MUX21_709 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n24), .Y(U[26]) );
  MUX21_708 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n24), .Y(U[27]) );
  MUX21_707 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n24), .Y(U[28]) );
  MUX21_706 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n24), .Y(U[29]) );
  MUX21_705 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n24), .Y(U[30]) );
  MUX21_704 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n24), .Y(U[31]) );
  BUF_X1 U1 ( .A(n21), .Z(n22) );
  BUF_X1 U2 ( .A(n21), .Z(n23) );
  BUF_X1 U3 ( .A(n21), .Z(n24) );
endmodule


module MUX21_40 ( in1, in0, S, Y );
  input in1, in0, S;
  output Y;
  wire   n3, n8;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(in0), .A2(n8), .B1(in1), .B2(S), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n8) );
endmodule


module mux21N_N32_16 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   n41, n42, n43, n44;
  assign n41 = S;

  MUX21_767 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n44), .Y(U[0]) );
  MUX21_766 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n42), .Y(U[1]) );
  MUX21_765 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n42), .Y(U[2]) );
  MUX21_764 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n42), .Y(U[3]) );
  MUX21_763 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n42), .Y(U[4]) );
  MUX21_762 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n42), .Y(U[5]) );
  MUX21_761 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n42), .Y(U[6]) );
  MUX21_760 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n42), .Y(U[7]) );
  MUX21_759 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n42), .Y(U[8]) );
  MUX21_758 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n42), .Y(U[9]) );
  MUX21_757 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n42), .Y(U[10]) );
  MUX21_756 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n42), .Y(U[11]) );
  MUX21_755 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n42), .Y(U[12]) );
  MUX21_754 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n43), .Y(U[13]) );
  MUX21_753 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n43), .Y(U[14]) );
  MUX21_752 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n43), .Y(U[15]) );
  MUX21_751 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n43), .Y(U[16]) );
  MUX21_750 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n43), .Y(U[17]) );
  MUX21_749 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n43), .Y(U[18]) );
  MUX21_748 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n43), .Y(U[19]) );
  MUX21_747 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n43), .Y(U[20]) );
  MUX21_746 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n43), .Y(U[21]) );
  MUX21_745 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n43), .Y(U[22]) );
  MUX21_744 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n43), .Y(U[23]) );
  MUX21_743 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n43), .Y(U[24]) );
  MUX21_742 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n44), .Y(U[25]) );
  MUX21_741 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n44), .Y(U[26]) );
  MUX21_740 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n44), .Y(U[27]) );
  MUX21_739 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n44), .Y(U[28]) );
  MUX21_738 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n44), .Y(U[29]) );
  MUX21_737 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n44), .Y(U[30]) );
  MUX21_736 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n44), .Y(U[31]) );
  BUF_X2 U1 ( .A(n41), .Z(n43) );
  BUF_X2 U2 ( .A(n41), .Z(n42) );
  BUF_X2 U3 ( .A(n41), .Z(n44) );
endmodule


module PC_RAM_DEPTH30 ( PC_In, En, Clk, Res, PC_DATAP, PC_IRAM );
  input [31:0] PC_In;
  output [31:0] PC_DATAP;
  output [29:0] PC_IRAM;
  input En, Clk, Res;
  wire   n112, n113, n114, n115, n116, n117, n118;

  DFFR_X1 \PC_IRAM_reg[29]  ( .D(PC_In[31]), .CK(Clk), .RN(n115), .Q(
        PC_IRAM[29]) );
  DFFR_X1 \PC_IRAM_reg[28]  ( .D(PC_In[30]), .CK(Clk), .RN(n114), .Q(
        PC_IRAM[28]) );
  DFFR_X1 \PC_IRAM_reg[27]  ( .D(PC_In[29]), .CK(Clk), .RN(n114), .Q(
        PC_IRAM[27]) );
  DFFR_X1 \PC_IRAM_reg[26]  ( .D(PC_In[28]), .CK(Clk), .RN(n114), .Q(
        PC_IRAM[26]) );
  DFFR_X1 \PC_IRAM_reg[25]  ( .D(PC_In[27]), .CK(Clk), .RN(n115), .Q(
        PC_IRAM[25]) );
  DFFR_X1 \PC_IRAM_reg[24]  ( .D(PC_In[26]), .CK(Clk), .RN(n114), .Q(
        PC_IRAM[24]) );
  DFFR_X1 \PC_IRAM_reg[23]  ( .D(PC_In[25]), .CK(Clk), .RN(n114), .Q(
        PC_IRAM[23]) );
  DFFR_X1 \PC_IRAM_reg[22]  ( .D(PC_In[24]), .CK(Clk), .RN(n112), .Q(
        PC_IRAM[22]) );
  DFFR_X1 \PC_IRAM_reg[21]  ( .D(PC_In[23]), .CK(Clk), .RN(n115), .Q(
        PC_IRAM[21]) );
  DFFR_X1 \PC_IRAM_reg[20]  ( .D(PC_In[22]), .CK(Clk), .RN(n112), .Q(
        PC_IRAM[20]) );
  DFFR_X1 \PC_IRAM_reg[19]  ( .D(PC_In[21]), .CK(Clk), .RN(n112), .Q(
        PC_IRAM[19]) );
  DFFR_X1 \PC_IRAM_reg[18]  ( .D(PC_In[20]), .CK(Clk), .RN(n112), .Q(
        PC_IRAM[18]) );
  DFFR_X1 \PC_IRAM_reg[17]  ( .D(PC_In[19]), .CK(Clk), .RN(n115), .Q(
        PC_IRAM[17]) );
  DFFR_X1 \PC_IRAM_reg[16]  ( .D(PC_In[18]), .CK(Clk), .RN(n112), .Q(
        PC_IRAM[16]) );
  DFFR_X1 \PC_IRAM_reg[15]  ( .D(PC_In[17]), .CK(Clk), .RN(n117), .Q(
        PC_IRAM[15]) );
  DFFR_X1 \PC_IRAM_reg[14]  ( .D(PC_In[16]), .CK(Clk), .RN(n113), .Q(
        PC_IRAM[14]) );
  DFFR_X1 \PC_IRAM_reg[13]  ( .D(PC_In[15]), .CK(Clk), .RN(n115), .Q(
        PC_IRAM[13]) );
  DFFR_X1 \PC_IRAM_reg[12]  ( .D(PC_In[14]), .CK(Clk), .RN(n113), .Q(
        PC_IRAM[12]) );
  DFFR_X1 \PC_IRAM_reg[11]  ( .D(PC_In[13]), .CK(Clk), .RN(n113), .Q(
        PC_IRAM[11]) );
  DFFR_X1 \PC_IRAM_reg[10]  ( .D(PC_In[12]), .CK(Clk), .RN(n113), .Q(
        PC_IRAM[10]) );
  DFFR_X1 \PC_IRAM_reg[9]  ( .D(PC_In[11]), .CK(Clk), .RN(n115), .Q(PC_IRAM[9]) );
  DFFR_X1 \PC_IRAM_reg[8]  ( .D(PC_In[10]), .CK(Clk), .RN(n113), .Q(PC_IRAM[8]) );
  DFFR_X1 \PC_IRAM_reg[7]  ( .D(PC_In[9]), .CK(Clk), .RN(n113), .Q(PC_IRAM[7])
         );
  DFFR_X1 \PC_IRAM_reg[6]  ( .D(PC_In[8]), .CK(Clk), .RN(n116), .Q(PC_IRAM[6])
         );
  DFFR_X1 \PC_IRAM_reg[5]  ( .D(PC_In[7]), .CK(Clk), .RN(n112), .Q(PC_IRAM[5])
         );
  DFFR_X1 \PC_IRAM_reg[4]  ( .D(PC_In[6]), .CK(Clk), .RN(n116), .Q(PC_IRAM[4])
         );
  DFFR_X1 \PC_IRAM_reg[3]  ( .D(PC_In[5]), .CK(Clk), .RN(n116), .Q(PC_IRAM[3])
         );
  DFFR_X1 \PC_IRAM_reg[2]  ( .D(PC_In[4]), .CK(Clk), .RN(n116), .Q(PC_IRAM[2])
         );
  DFFR_X1 \PC_IRAM_reg[1]  ( .D(PC_In[3]), .CK(Clk), .RN(n116), .Q(PC_IRAM[1])
         );
  DFFR_X1 \PC_IRAM_reg[0]  ( .D(PC_In[2]), .CK(Clk), .RN(n116), .Q(PC_IRAM[0])
         );
  DFFR_X1 \PC_DATAP_reg[31]  ( .D(PC_In[31]), .CK(Clk), .RN(n114), .Q(
        PC_DATAP[31]) );
  DFFR_X1 \PC_DATAP_reg[30]  ( .D(PC_In[30]), .CK(Clk), .RN(n114), .Q(
        PC_DATAP[30]) );
  DFFR_X1 \PC_DATAP_reg[29]  ( .D(PC_In[29]), .CK(Clk), .RN(n114), .Q(
        PC_DATAP[29]) );
  DFFR_X1 \PC_DATAP_reg[28]  ( .D(PC_In[28]), .CK(Clk), .RN(n114), .Q(
        PC_DATAP[28]) );
  DFFR_X1 \PC_DATAP_reg[27]  ( .D(PC_In[27]), .CK(Clk), .RN(n115), .Q(
        PC_DATAP[27]) );
  DFFR_X1 \PC_DATAP_reg[26]  ( .D(PC_In[26]), .CK(Clk), .RN(n114), .Q(
        PC_DATAP[26]) );
  DFFR_X1 \PC_DATAP_reg[25]  ( .D(PC_In[25]), .CK(Clk), .RN(n114), .Q(
        PC_DATAP[25]) );
  DFFR_X1 \PC_DATAP_reg[24]  ( .D(PC_In[24]), .CK(Clk), .RN(n114), .Q(
        PC_DATAP[24]) );
  DFFR_X1 \PC_DATAP_reg[23]  ( .D(PC_In[23]), .CK(Clk), .RN(n115), .Q(
        PC_DATAP[23]) );
  DFFR_X1 \PC_DATAP_reg[22]  ( .D(PC_In[22]), .CK(Clk), .RN(n112), .Q(
        PC_DATAP[22]) );
  DFFR_X1 \PC_DATAP_reg[21]  ( .D(PC_In[21]), .CK(Clk), .RN(n112), .Q(
        PC_DATAP[21]) );
  DFFR_X1 \PC_DATAP_reg[20]  ( .D(PC_In[20]), .CK(Clk), .RN(n112), .Q(
        PC_DATAP[20]) );
  DFFR_X1 \PC_DATAP_reg[19]  ( .D(PC_In[19]), .CK(Clk), .RN(n115), .Q(
        PC_DATAP[19]) );
  DFFR_X1 \PC_DATAP_reg[18]  ( .D(PC_In[18]), .CK(Clk), .RN(n112), .Q(
        PC_DATAP[18]) );
  DFFR_X1 \PC_DATAP_reg[17]  ( .D(PC_In[17]), .CK(Clk), .RN(n112), .Q(
        PC_DATAP[17]) );
  DFFR_X1 \PC_DATAP_reg[16]  ( .D(PC_In[16]), .CK(Clk), .RN(n117), .Q(
        PC_DATAP[16]) );
  DFFR_X1 \PC_DATAP_reg[15]  ( .D(PC_In[15]), .CK(Clk), .RN(n115), .Q(
        PC_DATAP[15]) );
  DFFR_X1 \PC_DATAP_reg[14]  ( .D(PC_In[14]), .CK(Clk), .RN(n113), .Q(
        PC_DATAP[14]) );
  DFFR_X1 \PC_DATAP_reg[13]  ( .D(PC_In[13]), .CK(Clk), .RN(n113), .Q(
        PC_DATAP[13]) );
  DFFR_X1 \PC_DATAP_reg[12]  ( .D(PC_In[12]), .CK(Clk), .RN(n113), .Q(
        PC_DATAP[12]) );
  DFFR_X1 \PC_DATAP_reg[11]  ( .D(PC_In[11]), .CK(Clk), .RN(n115), .Q(
        PC_DATAP[11]) );
  DFFR_X1 \PC_DATAP_reg[10]  ( .D(PC_In[10]), .CK(Clk), .RN(n113), .Q(
        PC_DATAP[10]) );
  DFFR_X1 \PC_DATAP_reg[9]  ( .D(PC_In[9]), .CK(Clk), .RN(n113), .Q(
        PC_DATAP[9]) );
  DFFR_X1 \PC_DATAP_reg[8]  ( .D(PC_In[8]), .CK(Clk), .RN(n113), .Q(
        PC_DATAP[8]) );
  DFFR_X1 \PC_DATAP_reg[7]  ( .D(PC_In[7]), .CK(Clk), .RN(n115), .Q(
        PC_DATAP[7]) );
  DFFR_X1 \PC_DATAP_reg[6]  ( .D(PC_In[6]), .CK(Clk), .RN(n116), .Q(
        PC_DATAP[6]) );
  DFFR_X1 \PC_DATAP_reg[5]  ( .D(PC_In[5]), .CK(Clk), .RN(n116), .Q(
        PC_DATAP[5]) );
  DFFR_X1 \PC_DATAP_reg[4]  ( .D(PC_In[4]), .CK(Clk), .RN(n116), .Q(
        PC_DATAP[4]) );
  DFFR_X1 \PC_DATAP_reg[3]  ( .D(PC_In[3]), .CK(Clk), .RN(n116), .Q(
        PC_DATAP[3]) );
  DFFR_X1 \PC_DATAP_reg[2]  ( .D(PC_In[2]), .CK(Clk), .RN(n116), .Q(
        PC_DATAP[2]) );
  DFFR_X1 \PC_DATAP_reg[1]  ( .D(PC_In[1]), .CK(Clk), .RN(n116), .Q(
        PC_DATAP[1]) );
  DFFR_X1 \PC_DATAP_reg[0]  ( .D(PC_In[0]), .CK(Clk), .RN(n112), .Q(
        PC_DATAP[0]) );
  CLKBUF_X1 U3 ( .A(n118), .Z(n112) );
  CLKBUF_X1 U4 ( .A(n118), .Z(n113) );
  CLKBUF_X1 U5 ( .A(n118), .Z(n114) );
  CLKBUF_X1 U6 ( .A(n118), .Z(n115) );
  CLKBUF_X1 U7 ( .A(n118), .Z(n116) );
  CLKBUF_X1 U8 ( .A(n118), .Z(n117) );
  INV_X1 U9 ( .A(Res), .ZN(n118) );
endmodule


module mux21N_N32_0 ( in1, in0, S, U );
  input [31:0] in1;
  input [31:0] in0;
  output [31:0] U;
  input S;
  wire   n24, n25, n26, n27;
  assign n24 = S;

  MUX21_799 muxes_0 ( .in1(in1[0]), .in0(in0[0]), .S(n27), .Y(U[0]) );
  MUX21_798 muxes_1 ( .in1(in1[1]), .in0(in0[1]), .S(n27), .Y(U[1]) );
  MUX21_797 muxes_2 ( .in1(in1[2]), .in0(in0[2]), .S(n27), .Y(U[2]) );
  MUX21_796 muxes_3 ( .in1(in1[3]), .in0(in0[3]), .S(n27), .Y(U[3]) );
  MUX21_795 muxes_4 ( .in1(in1[4]), .in0(in0[4]), .S(n27), .Y(U[4]) );
  MUX21_794 muxes_5 ( .in1(in1[5]), .in0(in0[5]), .S(n27), .Y(U[5]) );
  MUX21_793 muxes_6 ( .in1(in1[6]), .in0(in0[6]), .S(n27), .Y(U[6]) );
  MUX21_792 muxes_7 ( .in1(in1[7]), .in0(in0[7]), .S(n27), .Y(U[7]) );
  MUX21_791 muxes_8 ( .in1(in1[8]), .in0(in0[8]), .S(n25), .Y(U[8]) );
  MUX21_790 muxes_9 ( .in1(in1[9]), .in0(in0[9]), .S(n25), .Y(U[9]) );
  MUX21_789 muxes_10 ( .in1(in1[10]), .in0(in0[10]), .S(n25), .Y(U[10]) );
  MUX21_788 muxes_11 ( .in1(in1[11]), .in0(in0[11]), .S(n25), .Y(U[11]) );
  MUX21_787 muxes_12 ( .in1(in1[12]), .in0(in0[12]), .S(n25), .Y(U[12]) );
  MUX21_786 muxes_13 ( .in1(in1[13]), .in0(in0[13]), .S(n25), .Y(U[13]) );
  MUX21_785 muxes_14 ( .in1(in1[14]), .in0(in0[14]), .S(n25), .Y(U[14]) );
  MUX21_784 muxes_15 ( .in1(in1[15]), .in0(in0[15]), .S(n25), .Y(U[15]) );
  MUX21_783 muxes_16 ( .in1(in1[16]), .in0(in0[16]), .S(n25), .Y(U[16]) );
  MUX21_782 muxes_17 ( .in1(in1[17]), .in0(in0[17]), .S(n25), .Y(U[17]) );
  MUX21_781 muxes_18 ( .in1(in1[18]), .in0(in0[18]), .S(n25), .Y(U[18]) );
  MUX21_780 muxes_19 ( .in1(in1[19]), .in0(in0[19]), .S(n25), .Y(U[19]) );
  MUX21_779 muxes_20 ( .in1(in1[20]), .in0(in0[20]), .S(n26), .Y(U[20]) );
  MUX21_778 muxes_21 ( .in1(in1[21]), .in0(in0[21]), .S(n26), .Y(U[21]) );
  MUX21_777 muxes_22 ( .in1(in1[22]), .in0(in0[22]), .S(n26), .Y(U[22]) );
  MUX21_776 muxes_23 ( .in1(in1[23]), .in0(in0[23]), .S(n26), .Y(U[23]) );
  MUX21_775 muxes_24 ( .in1(in1[24]), .in0(in0[24]), .S(n26), .Y(U[24]) );
  MUX21_774 muxes_25 ( .in1(in1[25]), .in0(in0[25]), .S(n26), .Y(U[25]) );
  MUX21_773 muxes_26 ( .in1(in1[26]), .in0(in0[26]), .S(n26), .Y(U[26]) );
  MUX21_772 muxes_27 ( .in1(in1[27]), .in0(in0[27]), .S(n26), .Y(U[27]) );
  MUX21_771 muxes_28 ( .in1(in1[28]), .in0(in0[28]), .S(n26), .Y(U[28]) );
  MUX21_770 muxes_29 ( .in1(in1[29]), .in0(in0[29]), .S(n26), .Y(U[29]) );
  MUX21_769 muxes_30 ( .in1(in1[30]), .in0(in0[30]), .S(n26), .Y(U[30]) );
  MUX21_768 muxes_31 ( .in1(in1[31]), .in0(in0[31]), .S(n26), .Y(U[31]) );
  BUF_X1 U1 ( .A(n24), .Z(n25) );
  BUF_X1 U2 ( .A(n24), .Z(n26) );
  CLKBUF_X1 U3 ( .A(n24), .Z(n27) );
endmodule


module CU_HW_FUNC_SIZE11_OP_CODE_SIZE6_NALUop4_I_SIZE32_CW_SIZE42 ( Clk, Rst, 
        Inst, BrNZ, BrZ, BranchInst, StoreInst, JumpRInst, LHIInst, FS_Rst, 
        FATCHRstMux21_Sel, FATCH_En, PCMux41_Sel, Jump, IRAM_Rst, DECODE_Rst, 
        DECODE_En, RF_Rst, RF_RD1, RF_RD2, R1Mux21A_Sel, R2Mux21B_Sel, 
        RWMux41WR_Sel, ImmMux21_Sel, EXECUTE_Rst, EXECUTE_En, OPAMux21_Sel, 
        OPBMux41_Sel, ALU_Sel, ALU_Unsign, ALU_Arith_logN, StatusMux81_sel, 
        MEMORY_Rst, MEMORY_En, DATAMEM_En, DATAMEM_Rst, DATAMEM_Read_Wrn, 
        DATAMEM_Word, DATAMEM_HalfWord, DATAMEM_Byte, DATAMEM_Unsign, RF_WR, 
        WBMux41_Sel );
  input [31:0] Inst;
  output [1:0] PCMux41_Sel;
  output [1:0] RWMux41WR_Sel;
  output [1:0] OPBMux41_Sel;
  output [3:0] ALU_Sel;
  output [2:0] StatusMux81_sel;
  output [1:0] WBMux41_Sel;
  input Clk, Rst, BrNZ, BrZ;
  output BranchInst, StoreInst, JumpRInst, LHIInst, FS_Rst, FATCHRstMux21_Sel,
         FATCH_En, Jump, IRAM_Rst, DECODE_Rst, DECODE_En, RF_Rst, RF_RD1,
         RF_RD2, R1Mux21A_Sel, R2Mux21B_Sel, ImmMux21_Sel, EXECUTE_Rst,
         EXECUTE_En, OPAMux21_Sel, ALU_Unsign, ALU_Arith_logN, MEMORY_Rst,
         MEMORY_En, DATAMEM_En, DATAMEM_Rst, DATAMEM_Read_Wrn, DATAMEM_Word,
         DATAMEM_HalfWord, DATAMEM_Byte, DATAMEM_Unsign, RF_WR;
  wire   Inst_31, Inst_30, Inst_29, Inst_28, Inst_27, Inst_26, notClk, N3792,
         N3793, N3794, n199, n202, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n234,
         n235, n236, n237, n238, n239, n240, n242, n244, n245, n246, n248,
         n250, n252, n254, n257, n260, n263, n266, n269, n273, n277, n281,
         n285, n289, n293, n297, n302, n307, n312, n317, n323, n329, n335,
         n340, n345, n350, n355, n360, n364, n368, n372, n376, n380, n384,
         n388, n391, n394, n397, n400, n403, n405, n407, n409, n413, n415,
         n417, n419, n421, n423, n425, n427, n429, n431, n433, n435, n437,
         n439, n441, n443, n445, n447, n449, n451, n453, n455, n457, n459,
         n461, n463, n465, n467, n469, n471, n473, n475, n477, n479, n481,
         n483, n485, n487, n489, n491, n493, n495, n497, n499, n501, n503,
         n505, n507, n509, n511, n513, n515, n517, n519, n521, n523, n525,
         n527, n529, n531, n533, n535, n537, n539, n541, n543, n545, n547,
         n549, n551, n553, n555, n557, n559, n561, n563, n565, n567, n569,
         n571, n573, n575, n577, n579, n581, n583, n585, n587, n589, n591,
         n593, n595, n597, n599, n601, n603, n605, n607, n609, n611, n613,
         n615, n617, n620, n622, n624, n626, n628, n630, n632, n634, n636,
         n639, n642, n643, n295, n280, n709, n711, n48, n49, n50, n52, n53,
         n54, n55, n56, n57, n58, n59, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n183, n184, n185, n187,
         n188, n189, n191, n192, n193, n194, n195, n196, n197, n198, n200,
         n215, n233, n241, n243, n249, n251, n253, n255, n256, n258, n259,
         n261, n262, n264, n265, n267, n268, n270, n271, n272, n274, n275,
         n276, n278, n279, n282, n283, n751, n752, n753, n754, n759, n761,
         n763, n765, n767, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783;
  wire   [41:0] CW;
  tri   FS_Rst;
  tri   FATCHRstMux21_Sel;
  tri   [1:0] PCMux41_Sel;
  tri   IRAM_Rst;
  tri   RF_Rst;
  tri   RF_RD1;
  tri   RF_RD2;
  tri   R1Mux21A_Sel;
  tri   R2Mux21B_Sel;
  tri   [1:0] RWMux41WR_Sel;
  tri   ImmMux21_Sel;
  tri   OPAMux21_Sel;
  tri   [1:0] OPBMux41_Sel;
  tri   [3:0] ALU_Sel;
  tri   ALU_Unsign;
  tri   ALU_Arith_logN;
  tri   [2:0] StatusMux81_sel;
  tri   DATAMEM_En;
  tri   DATAMEM_Rst;
  tri   DATAMEM_Read_Wrn;
  tri   DATAMEM_Word;
  tri   DATAMEM_HalfWord;
  tri   DATAMEM_Byte;
  tri   DATAMEM_Unsign;
  tri   RF_WR;
  tri   [35:0] CWSF;
  tri   [25:0] CWSD;
  tri   [11:0] CWSE;
  tri   [2:0] CWSM;
  tri   n784;
  tri   n791;
  tri   n789;
  tri   n787;
  tri   n792;
  tri   n788;
  tri   n790;
  tri   n785;
  tri   n786;
  assign Inst_31 = Inst[31];
  assign Inst_30 = Inst[30];
  assign Inst_29 = Inst[29];
  assign Inst_28 = Inst[28];
  assign Inst_27 = Inst[27];
  assign Inst_26 = Inst[26];

  DFF_X1 BranchNZ_In_reg ( .D(n643), .CK(Clk), .Q(n280), .QN(n709) );
  DFF_X1 \CW_reg[41]  ( .D(n642), .CK(Clk), .Q(CW[41]), .QN(n239) );
  DFF_X1 \CWSF_reg[41]  ( .D(CW[41]), .CK(notClk), .Q(FS_Rst) );
  DFF_X1 \CW_reg[39]  ( .D(n639), .CK(Clk), .Q(CW[39]), .QN(n238) );
  DFF_X1 \CWSF_reg[39]  ( .D(CW[39]), .CK(notClk), .Q(FATCHRstMux21_Sel) );
  DFF_X1 \CWSF_reg[36]  ( .D(1'b0), .CK(notClk), .Q(IRAM_Rst) );
  DFF_X1 \CW_reg[35]  ( .D(n636), .CK(Clk), .Q(CW[35]), .QN(n237) );
  DFF_X1 \CWSF_reg[35]  ( .D(CW[35]), .CK(notClk), .Q(CWSF[35]) );
  DFF_X1 \CW_reg[34]  ( .D(n634), .CK(Clk), .Q(CW[34]), .QN(n236) );
  DFF_X1 \CWSF_reg[34]  ( .D(CW[34]), .CK(notClk), .Q(CWSF[34]) );
  DFF_X1 \CW_reg[33]  ( .D(n632), .CK(Clk), .Q(CW[33]), .QN(n235) );
  DFF_X1 \CWSF_reg[33]  ( .D(CW[33]), .CK(notClk), .Q(CWSF[33]) );
  DFF_X1 \CW_reg[32]  ( .D(n630), .CK(Clk), .Q(CW[32]), .QN(n234) );
  DFF_X1 \CWSF_reg[32]  ( .D(CW[32]), .CK(notClk), .Q(CWSF[32]) );
  DFF_X1 \CW_reg[31]  ( .D(n628), .CK(Clk), .Q(CW[31]) );
  DFF_X1 \CWSF_reg[31]  ( .D(CW[31]), .CK(notClk), .Q(CWSF[31]) );
  DFF_X1 \CW_reg[30]  ( .D(n626), .CK(Clk), .Q(CW[30]), .QN(n232) );
  DFF_X1 \CWSF_reg[30]  ( .D(CW[30]), .CK(notClk), .Q(CWSF[30]) );
  DFF_X1 \CW_reg[29]  ( .D(n624), .CK(Clk), .Q(CW[29]), .QN(n231) );
  DFF_X1 \CWSF_reg[29]  ( .D(CW[29]), .CK(notClk), .Q(CWSF[29]) );
  DFF_X1 \CW_reg[28]  ( .D(n622), .CK(Clk), .Q(CW[28]), .QN(n230) );
  DFF_X1 \CWSF_reg[28]  ( .D(CW[28]), .CK(notClk), .Q(CWSF[28]) );
  DFF_X1 \CW_reg[27]  ( .D(n620), .CK(Clk), .Q(CW[27]), .QN(n229) );
  DFF_X1 \CWSF_reg[27]  ( .D(CW[27]), .CK(notClk), .Q(CWSF[27]) );
  DFF_X1 \CWSF_reg[26]  ( .D(1'b0), .CK(notClk), .Q(CWSF[26]) );
  DFF_X1 \CW_reg[25]  ( .D(n617), .CK(Clk), .Q(CW[25]), .QN(n228) );
  DFF_X1 \CWSF_reg[25]  ( .D(CW[25]), .CK(notClk), .Q(CWSF[25]) );
  DFF_X1 \CW_reg[24]  ( .D(n615), .CK(Clk), .Q(CW[24]), .QN(n227) );
  DFF_X1 \CWSF_reg[24]  ( .D(CW[24]), .CK(notClk), .Q(CWSF[24]) );
  DFF_X1 \CW_reg[23]  ( .D(n613), .CK(Clk), .Q(CW[23]), .QN(n226) );
  DFF_X1 \CWSF_reg[23]  ( .D(CW[23]), .CK(notClk), .Q(CWSF[23]) );
  DFF_X1 \CW_reg[22]  ( .D(n611), .CK(Clk), .Q(CW[22]), .QN(n225) );
  DFF_X1 \CWSF_reg[22]  ( .D(CW[22]), .CK(notClk), .Q(CWSF[22]) );
  DFF_X1 \CW_reg[21]  ( .D(n609), .CK(Clk), .Q(CW[21]), .QN(n224) );
  DFF_X1 \CWSF_reg[21]  ( .D(CW[21]), .CK(notClk), .Q(CWSF[21]) );
  DFF_X1 \CW_reg[20]  ( .D(n607), .CK(Clk), .Q(CW[20]), .QN(n223) );
  DFF_X1 \CWSF_reg[20]  ( .D(CW[20]), .CK(notClk), .Q(CWSF[20]) );
  DFF_X1 \CW_reg[19]  ( .D(n605), .CK(Clk), .Q(CW[19]), .QN(n222) );
  DFF_X1 \CWSF_reg[19]  ( .D(CW[19]), .CK(notClk), .Q(CWSF[19]) );
  DFF_X1 \CW_reg[18]  ( .D(n603), .CK(Clk), .Q(CW[18]), .QN(n221) );
  DFF_X1 \CWSF_reg[18]  ( .D(CW[18]), .CK(notClk), .Q(CWSF[18]) );
  DFF_X1 \CW_reg[17]  ( .D(n601), .CK(Clk), .Q(CW[17]), .QN(n220) );
  DFF_X1 \CWSF_reg[17]  ( .D(CW[17]), .CK(notClk), .Q(CWSF[17]) );
  DFF_X1 \CW_reg[16]  ( .D(n599), .CK(Clk), .Q(CW[16]), .QN(n219) );
  DFF_X1 \CWSF_reg[16]  ( .D(CW[16]), .CK(notClk), .Q(CWSF[16]) );
  DFF_X1 \CW_reg[15]  ( .D(n597), .CK(Clk), .Q(CW[15]), .QN(n218) );
  DFF_X1 \CWSF_reg[15]  ( .D(CW[15]), .CK(notClk), .Q(CWSF[15]) );
  DFF_X1 \CW_reg[14]  ( .D(n595), .CK(Clk), .Q(CW[14]), .QN(n217) );
  DFF_X1 \CWSF_reg[14]  ( .D(CW[14]), .CK(notClk), .Q(CWSF[14]) );
  DFF_X1 \CW_reg[13]  ( .D(n593), .CK(Clk), .Q(CW[13]), .QN(n216) );
  DFF_X1 \CWSF_reg[13]  ( .D(CW[13]), .CK(notClk), .Q(CWSF[13]) );
  DFF_X1 \CW_reg[12]  ( .D(n591), .CK(Clk), .Q(CW[12]), .QN(n295) );
  DFF_X1 \CWSF_reg[12]  ( .D(CW[12]), .CK(notClk), .Q(CWSF[12]) );
  DFF_X1 \CW_reg[11]  ( .D(n589), .CK(Clk), .Q(CW[11]), .QN(n214) );
  DFF_X1 \CWSF_reg[11]  ( .D(CW[11]), .CK(notClk), .Q(CWSF[11]) );
  DFF_X1 \CW_reg[10]  ( .D(n587), .CK(Clk), .Q(CW[10]), .QN(n213) );
  DFF_X1 \CWSF_reg[10]  ( .D(CW[10]), .CK(notClk), .Q(CWSF[10]) );
  DFF_X1 \CW_reg[9]  ( .D(n585), .CK(Clk), .Q(CW[9]), .QN(n212) );
  DFF_X1 \CWSF_reg[9]  ( .D(CW[9]), .CK(notClk), .Q(CWSF[9]) );
  DFF_X1 \CW_reg[8]  ( .D(n583), .CK(Clk), .Q(CW[8]), .QN(n211) );
  DFF_X1 \CWSF_reg[8]  ( .D(CW[8]), .CK(notClk), .Q(CWSF[8]) );
  DFF_X1 \CW_reg[7]  ( .D(n581), .CK(Clk), .Q(CW[7]), .QN(n210) );
  DFF_X1 \CWSF_reg[7]  ( .D(CW[7]), .CK(notClk), .Q(CWSF[7]) );
  DFF_X1 \CW_reg[6]  ( .D(n579), .CK(Clk), .Q(CW[6]), .QN(n209) );
  DFF_X1 \CWSF_reg[6]  ( .D(CW[6]), .CK(notClk), .Q(CWSF[6]) );
  DFF_X1 \CW_reg[5]  ( .D(n577), .CK(Clk), .Q(CW[5]), .QN(n208) );
  DFF_X1 \CWSF_reg[5]  ( .D(CW[5]), .CK(notClk), .Q(CWSF[5]) );
  DFF_X1 \CW_reg[4]  ( .D(n575), .CK(Clk), .Q(CW[4]), .QN(n207) );
  DFF_X1 \CWSF_reg[4]  ( .D(CW[4]), .CK(notClk), .Q(CWSF[4]) );
  DFF_X1 \CW_reg[3]  ( .D(n573), .CK(Clk), .Q(CW[3]), .QN(n206) );
  DFF_X1 \CWSF_reg[3]  ( .D(CW[3]), .CK(notClk), .Q(CWSF[3]) );
  DFF_X1 \CW_reg[2]  ( .D(n571), .CK(Clk), .Q(CW[2]), .QN(n205) );
  DFF_X1 \CWSF_reg[2]  ( .D(CW[2]), .CK(notClk), .Q(CWSF[2]) );
  DFF_X1 \CW_reg[1]  ( .D(n569), .CK(Clk), .Q(CW[1]), .QN(n204) );
  DFF_X1 \CWSF_reg[1]  ( .D(CW[1]), .CK(notClk), .Q(CWSF[1]) );
  DFF_X1 \CW_reg[0]  ( .D(n567), .CK(Clk), .Q(CW[0]) );
  DFF_X1 \CWSF_reg[0]  ( .D(CW[0]), .CK(notClk), .Q(CWSF[0]) );
  DFF_X1 \CWSD_reg2[35]  ( .D(n565), .CK(Clk), .Q(n786) );
  DFF_X1 \CWSD_reg2[34]  ( .D(n563), .CK(Clk), .Q(n785) );
  DFF_X1 \CWSD_reg2[33]  ( .D(n561), .CK(Clk), .Q(RF_Rst) );
  DFF_X1 \CWSD_reg2[32]  ( .D(n559), .CK(Clk), .Q(RF_RD1) );
  DFF_X1 \CWSD_reg2[31]  ( .D(n557), .CK(Clk), .Q(RF_RD2) );
  DFF_X1 \CWSD_reg2[30]  ( .D(n555), .CK(Clk), .Q(R1Mux21A_Sel) );
  DFF_X1 \CWSD_reg2[29]  ( .D(n553), .CK(Clk), .Q(R2Mux21B_Sel) );
  DFF_X1 \CWSD_reg2[28]  ( .D(n551), .CK(Clk), .Q(RWMux41WR_Sel[1]) );
  DFF_X1 \CWSD_reg2[27]  ( .D(n549), .CK(Clk), .Q(RWMux41WR_Sel[0]) );
  DFF_X1 \CWSD_reg2[26]  ( .D(n547), .CK(Clk), .Q(ImmMux21_Sel) );
  DFF_X1 \CWSD_reg2[25]  ( .D(n545), .CK(Clk), .Q(CWSD[25]) );
  DFF_X1 \CWSD_reg2[24]  ( .D(n543), .CK(Clk), .Q(CWSD[24]) );
  DFF_X1 \CWSD_reg2[23]  ( .D(n541), .CK(Clk), .Q(CWSD[23]) );
  DFF_X1 \CWSD_reg2[22]  ( .D(n539), .CK(Clk), .Q(CWSD[22]) );
  DFF_X1 \CWSD_reg2[21]  ( .D(n537), .CK(Clk), .Q(CWSD[21]) );
  DFF_X1 \CWSD_reg2[20]  ( .D(n535), .CK(Clk), .Q(CWSD[20]) );
  DFF_X1 \CWSD_reg2[19]  ( .D(n533), .CK(Clk), .Q(CWSD[19]) );
  DFF_X1 \CWSD_reg2[18]  ( .D(n531), .CK(Clk), .Q(CWSD[18]) );
  DFF_X1 \CWSD_reg2[17]  ( .D(n529), .CK(Clk), .Q(CWSD[17]) );
  DFF_X1 \CWSD_reg2[16]  ( .D(n527), .CK(Clk), .Q(CWSD[16]) );
  DFF_X1 \CWSD_reg2[15]  ( .D(n525), .CK(Clk), .Q(CWSD[15]) );
  DFF_X1 \CWSD_reg2[14]  ( .D(n523), .CK(Clk), .Q(CWSD[14]) );
  DFF_X1 \CWSD_reg2[13]  ( .D(n521), .CK(Clk), .Q(CWSD[13]) );
  DFF_X1 \CWSD_reg2[12]  ( .D(n519), .CK(Clk), .Q(CWSD[12]) );
  DFF_X1 \CWSD_reg2[11]  ( .D(n517), .CK(Clk), .Q(CWSD[11]) );
  DFF_X1 \CWSD_reg2[10]  ( .D(n515), .CK(Clk), .Q(CWSD[10]) );
  DFF_X1 \CWSD_reg2[9]  ( .D(n513), .CK(Clk), .Q(CWSD[9]) );
  DFF_X1 \CWSD_reg2[8]  ( .D(n511), .CK(Clk), .Q(CWSD[8]) );
  DFF_X1 \CWSD_reg2[7]  ( .D(n509), .CK(Clk), .Q(CWSD[7]) );
  DFF_X1 \CWSD_reg2[6]  ( .D(n507), .CK(Clk), .Q(CWSD[6]) );
  DFF_X1 \CWSD_reg2[5]  ( .D(n505), .CK(Clk), .Q(CWSD[5]) );
  DFF_X1 \CWSD_reg2[4]  ( .D(n503), .CK(Clk), .Q(CWSD[4]) );
  DFF_X1 \CWSD_reg2[3]  ( .D(n501), .CK(Clk), .Q(CWSD[3]) );
  DFF_X1 \CWSD_reg2[2]  ( .D(n499), .CK(Clk), .Q(CWSD[2]) );
  DFF_X1 \CWSD_reg2[1]  ( .D(n497), .CK(Clk), .Q(CWSD[1]) );
  DFF_X1 \CWSD_reg2[0]  ( .D(n495), .CK(Clk), .Q(CWSD[0]) );
  DFF_X1 \CWSE_reg2[25]  ( .D(n493), .CK(Clk), .Q(n788) );
  DFF_X1 \CWSE_reg2[24]  ( .D(n491), .CK(Clk), .Q(n787) );
  DFF_X1 \CWSE_reg2[20]  ( .D(n483), .CK(Clk), .Q(ALU_Sel[3]) );
  DFF_X1 \CWSE_reg2[19]  ( .D(n481), .CK(Clk), .Q(ALU_Sel[2]) );
  DFF_X1 \CWSE_reg2[18]  ( .D(n479), .CK(Clk), .Q(ALU_Sel[1]) );
  DFF_X1 \CWSE_reg2[17]  ( .D(n477), .CK(Clk), .Q(ALU_Sel[0]) );
  DFF_X1 \CWSE_reg2[16]  ( .D(n475), .CK(Clk), .Q(ALU_Unsign) );
  DFF_X1 \CWSE_reg2[15]  ( .D(n473), .CK(Clk), .Q(ALU_Arith_logN) );
  DFF_X1 \CWSE_reg2[14]  ( .D(n471), .CK(Clk), .Q(StatusMux81_sel[2]) );
  DFF_X1 \CWSE_reg2[13]  ( .D(n469), .CK(Clk), .Q(StatusMux81_sel[1]) );
  DFF_X1 \CWSE_reg2[12]  ( .D(n467), .CK(Clk), .Q(StatusMux81_sel[0]) );
  DFF_X1 \CWSE_reg2[11]  ( .D(n465), .CK(Clk), .Q(CWSE[11]) );
  DFF_X1 \CWSE_reg2[10]  ( .D(n463), .CK(Clk), .Q(CWSE[10]) );
  DFF_X1 \CWSE_reg2[9]  ( .D(n461), .CK(Clk), .Q(CWSE[9]) );
  DFF_X1 \CWSE_reg2[8]  ( .D(n459), .CK(Clk), .Q(CWSE[8]) );
  DFF_X1 \CWSE_reg2[7]  ( .D(n457), .CK(Clk), .Q(CWSE[7]) );
  DFF_X1 \CWSE_reg2[6]  ( .D(n455), .CK(Clk), .Q(CWSE[6]) );
  DFF_X1 \CWSE_reg2[5]  ( .D(n453), .CK(Clk), .Q(CWSE[5]) );
  DFF_X1 \CWSE_reg2[4]  ( .D(n451), .CK(Clk), .Q(CWSE[4]) );
  DFF_X1 \CWSE_reg2[3]  ( .D(n449), .CK(Clk), .Q(CWSE[3]) );
  DFF_X1 \CWSE_reg2[2]  ( .D(n447), .CK(Clk), .Q(CWSE[2]) );
  DFF_X1 \CWSE_reg2[1]  ( .D(n445), .CK(Clk), .Q(CWSE[1]) );
  DFF_X1 \CWSE_reg2[0]  ( .D(n443), .CK(Clk), .Q(CWSE[0]) );
  DFF_X1 \CWSM_reg2[11]  ( .D(n441), .CK(Clk), .Q(n790) );
  DFF_X1 \CWSM_reg2[10]  ( .D(n439), .CK(Clk), .Q(n789) );
  DFF_X1 \CWSM_reg2[9]  ( .D(n437), .CK(Clk), .Q(DATAMEM_En) );
  DFF_X1 \CWSM_reg2[8]  ( .D(n435), .CK(Clk), .Q(DATAMEM_Rst) );
  DFF_X1 \CWSM_reg2[7]  ( .D(n433), .CK(Clk), .Q(DATAMEM_Read_Wrn) );
  DFF_X1 \CWSM_reg2[6]  ( .D(n431), .CK(Clk), .Q(DATAMEM_Word) );
  DFF_X1 \CWSM_reg2[5]  ( .D(n429), .CK(Clk), .Q(DATAMEM_HalfWord) );
  DFF_X1 \CWSM_reg2[4]  ( .D(n427), .CK(Clk), .Q(DATAMEM_Byte) );
  DFF_X1 \CWSM_reg2[3]  ( .D(n425), .CK(Clk), .Q(DATAMEM_Unsign) );
  DFF_X1 \CWSM_reg2[2]  ( .D(n423), .CK(Clk), .Q(CWSM[2]) );
  DFF_X1 \CWSM_reg2[1]  ( .D(n421), .CK(Clk), .Q(CWSM[1]) );
  DFF_X1 \CWSM_reg2[0]  ( .D(n419), .CK(Clk), .Q(CWSM[0]) );
  DFF_X1 \CWSWB_reg2[2]  ( .D(n417), .CK(Clk), .Q(RF_WR) );
  DFF_X1 \CWSWB_reg2[1]  ( .D(n415), .CK(Clk), .Q(n791) );
  DFF_X1 \CWSWB_reg2[0]  ( .D(n413), .CK(Clk), .Q(n792) );
  DFF_X1 StoreInst_reg ( .D(N3793), .CK(Clk), .Q(StoreInst) );
  DFF_X1 \CWSF_reg2[41]  ( .D(n409), .CK(Clk), .Q(FS_Rst) );
  DFF_X1 \CWSF_reg2[39]  ( .D(n407), .CK(Clk), .Q(FATCHRstMux21_Sel) );
  DFF_X1 \CWSF_reg2[37]  ( .D(n405), .CK(Clk), .Q(PCMux41_Sel[0]) );
  DFF_X1 \CWSF_reg2[35]  ( .D(n403), .CK(Clk), .Q(CWSF[35]) );
  DFF_X1 \CWSF_reg2[33]  ( .D(n400), .CK(Clk), .Q(CWSF[33]) );
  DFF_X1 \CWSD_reg[33]  ( .D(CWSF[33]), .CK(notClk), .Q(RF_Rst) );
  DFF_X1 \CWSF_reg2[31]  ( .D(n397), .CK(Clk), .Q(CWSF[31]) );
  DFF_X1 \CWSD_reg[31]  ( .D(CWSF[31]), .CK(notClk), .Q(RF_RD2) );
  DFF_X1 \CWSF_reg2[29]  ( .D(n394), .CK(Clk), .Q(CWSF[29]) );
  DFF_X1 \CWSD_reg[29]  ( .D(CWSF[29]), .CK(notClk), .Q(R2Mux21B_Sel) );
  DFF_X1 \CWSF_reg2[27]  ( .D(n391), .CK(Clk), .Q(CWSF[27]) );
  DFF_X1 \CWSD_reg[27]  ( .D(CWSF[27]), .CK(notClk), .Q(RWMux41WR_Sel[0]) );
  DFF_X1 \CWSF_reg2[25]  ( .D(n388), .CK(Clk), .Q(CWSF[25]) );
  DFF_X1 \CWSD_reg[25]  ( .D(CWSF[25]), .CK(notClk), .Q(CWSD[25]) );
  DFF_X1 \CWSF_reg2[23]  ( .D(n384), .CK(Clk), .Q(CWSF[23]) );
  DFF_X1 \CWSD_reg[23]  ( .D(CWSF[23]), .CK(notClk), .Q(CWSD[23]) );
  DFF_X1 \CWSF_reg2[21]  ( .D(n380), .CK(Clk), .Q(CWSF[21]) );
  DFF_X1 \CWSD_reg[21]  ( .D(CWSF[21]), .CK(notClk), .Q(CWSD[21]) );
  DFF_X1 \CWSF_reg2[19]  ( .D(n376), .CK(Clk), .Q(CWSF[19]) );
  DFF_X1 \CWSD_reg[19]  ( .D(CWSF[19]), .CK(notClk), .Q(CWSD[19]) );
  DFF_X1 \CWSE_reg[19]  ( .D(CWSD[19]), .CK(notClk), .Q(ALU_Sel[2]) );
  DFF_X1 \CWSF_reg2[17]  ( .D(n372), .CK(Clk), .Q(CWSF[17]) );
  DFF_X1 \CWSD_reg[17]  ( .D(CWSF[17]), .CK(notClk), .Q(CWSD[17]) );
  DFF_X1 \CWSE_reg[17]  ( .D(CWSD[17]), .CK(notClk), .Q(ALU_Sel[0]) );
  DFF_X1 \CWSF_reg2[15]  ( .D(n368), .CK(Clk), .Q(CWSF[15]) );
  DFF_X1 \CWSD_reg[15]  ( .D(CWSF[15]), .CK(notClk), .Q(CWSD[15]) );
  DFF_X1 \CWSE_reg[15]  ( .D(CWSD[15]), .CK(notClk), .Q(ALU_Arith_logN) );
  DFF_X1 \CWSF_reg2[13]  ( .D(n364), .CK(Clk), .Q(CWSF[13]) );
  DFF_X1 \CWSD_reg[13]  ( .D(CWSF[13]), .CK(notClk), .Q(CWSD[13]) );
  DFF_X1 \CWSE_reg[13]  ( .D(CWSD[13]), .CK(notClk), .Q(StatusMux81_sel[1]) );
  DFF_X1 \CWSF_reg2[11]  ( .D(n360), .CK(Clk), .Q(CWSF[11]) );
  DFF_X1 \CWSD_reg[11]  ( .D(CWSF[11]), .CK(notClk), .Q(CWSD[11]) );
  DFF_X1 \CWSE_reg[11]  ( .D(CWSD[11]), .CK(notClk), .Q(CWSE[11]) );
  DFF_X1 \CWSF_reg2[9]  ( .D(n355), .CK(Clk), .Q(CWSF[9]) );
  DFF_X1 \CWSD_reg[9]  ( .D(CWSF[9]), .CK(notClk), .Q(CWSD[9]) );
  DFF_X1 \CWSE_reg[9]  ( .D(CWSD[9]), .CK(notClk), .Q(CWSE[9]) );
  DFF_X1 \CWSM_reg[9]  ( .D(CWSE[9]), .CK(notClk), .Q(DATAMEM_En) );
  DFF_X1 \CWSF_reg2[7]  ( .D(n350), .CK(Clk), .Q(CWSF[7]) );
  DFF_X1 \CWSD_reg[7]  ( .D(CWSF[7]), .CK(notClk), .Q(CWSD[7]) );
  DFF_X1 \CWSE_reg[7]  ( .D(CWSD[7]), .CK(notClk), .Q(CWSE[7]) );
  DFF_X1 \CWSM_reg[7]  ( .D(CWSE[7]), .CK(notClk), .Q(DATAMEM_Read_Wrn) );
  DFF_X1 \CWSF_reg2[5]  ( .D(n345), .CK(Clk), .Q(CWSF[5]) );
  DFF_X1 \CWSD_reg[5]  ( .D(CWSF[5]), .CK(notClk), .Q(CWSD[5]) );
  DFF_X1 \CWSE_reg[5]  ( .D(CWSD[5]), .CK(notClk), .Q(CWSE[5]) );
  DFF_X1 \CWSM_reg[5]  ( .D(CWSE[5]), .CK(notClk), .Q(DATAMEM_HalfWord) );
  DFF_X1 \CWSF_reg2[3]  ( .D(n340), .CK(Clk), .Q(CWSF[3]) );
  DFF_X1 \CWSD_reg[3]  ( .D(CWSF[3]), .CK(notClk), .Q(CWSD[3]) );
  DFF_X1 \CWSE_reg[3]  ( .D(CWSD[3]), .CK(notClk), .Q(CWSE[3]) );
  DFF_X1 \CWSM_reg[3]  ( .D(CWSE[3]), .CK(notClk), .Q(DATAMEM_Unsign) );
  DFF_X1 \CWSF_reg2[1]  ( .D(n335), .CK(Clk), .Q(CWSF[1]) );
  DFF_X1 \CWSD_reg[1]  ( .D(CWSF[1]), .CK(notClk), .Q(CWSD[1]) );
  DFF_X1 \CWSE_reg[1]  ( .D(CWSD[1]), .CK(notClk), .Q(CWSE[1]) );
  DFF_X1 \CWSM_reg[1]  ( .D(CWSE[1]), .CK(notClk), .Q(CWSM[1]) );
  DFF_X1 \CWSWB_reg[1]  ( .D(CWSM[1]), .CK(notClk), .Q(n791) );
  DFF_X1 \CWSF_reg2[0]  ( .D(n329), .CK(Clk), .Q(CWSF[0]) );
  DFF_X1 \CWSD_reg[0]  ( .D(CWSF[0]), .CK(notClk), .Q(CWSD[0]) );
  DFF_X1 \CWSE_reg[0]  ( .D(CWSD[0]), .CK(notClk), .Q(CWSE[0]) );
  DFF_X1 \CWSM_reg[0]  ( .D(CWSE[0]), .CK(notClk), .Q(CWSM[0]) );
  DFF_X1 \CWSF_reg2[2]  ( .D(n323), .CK(Clk), .Q(CWSF[2]) );
  DFF_X1 \CWSD_reg[2]  ( .D(CWSF[2]), .CK(notClk), .Q(CWSD[2]) );
  DFF_X1 \CWSE_reg[2]  ( .D(CWSD[2]), .CK(notClk), .Q(CWSE[2]) );
  DFF_X1 \CWSM_reg[2]  ( .D(CWSE[2]), .CK(notClk), .Q(CWSM[2]) );
  DFF_X1 \CWSWB_reg[2]  ( .D(CWSM[2]), .CK(notClk), .Q(RF_WR) );
  DFF_X1 \CWSF_reg2[4]  ( .D(n317), .CK(Clk), .Q(CWSF[4]) );
  DFF_X1 \CWSD_reg[4]  ( .D(CWSF[4]), .CK(notClk), .Q(CWSD[4]) );
  DFF_X1 \CWSE_reg[4]  ( .D(CWSD[4]), .CK(notClk), .Q(CWSE[4]) );
  DFF_X1 \CWSM_reg[4]  ( .D(CWSE[4]), .CK(notClk), .Q(DATAMEM_Byte) );
  DFF_X1 \CWSF_reg2[6]  ( .D(n312), .CK(Clk), .Q(CWSF[6]) );
  DFF_X1 \CWSD_reg[6]  ( .D(CWSF[6]), .CK(notClk), .Q(CWSD[6]) );
  DFF_X1 \CWSE_reg[6]  ( .D(CWSD[6]), .CK(notClk), .Q(CWSE[6]) );
  DFF_X1 \CWSM_reg[6]  ( .D(CWSE[6]), .CK(notClk), .Q(DATAMEM_Word) );
  DFF_X1 \CWSF_reg2[8]  ( .D(n307), .CK(Clk), .Q(CWSF[8]) );
  DFF_X1 \CWSD_reg[8]  ( .D(CWSF[8]), .CK(notClk), .Q(CWSD[8]) );
  DFF_X1 \CWSE_reg[8]  ( .D(CWSD[8]), .CK(notClk), .Q(CWSE[8]) );
  DFF_X1 \CWSM_reg[8]  ( .D(CWSE[8]), .CK(notClk), .Q(DATAMEM_Rst) );
  DFF_X1 \CWSF_reg2[10]  ( .D(n302), .CK(Clk), .Q(CWSF[10]) );
  DFF_X1 \CWSD_reg[10]  ( .D(CWSF[10]), .CK(notClk), .Q(CWSD[10]) );
  DFF_X1 \CWSE_reg[10]  ( .D(CWSD[10]), .CK(notClk), .Q(CWSE[10]) );
  DFF_X1 \CWSF_reg2[12]  ( .D(n297), .CK(Clk), .Q(CWSF[12]) );
  DFF_X1 \CWSD_reg[12]  ( .D(CWSF[12]), .CK(notClk), .Q(CWSD[12]) );
  DFF_X1 \CWSE_reg[12]  ( .D(CWSD[12]), .CK(notClk), .Q(StatusMux81_sel[0]) );
  DFF_X1 \CWSF_reg2[14]  ( .D(n293), .CK(Clk), .Q(CWSF[14]) );
  DFF_X1 \CWSD_reg[14]  ( .D(CWSF[14]), .CK(notClk), .Q(CWSD[14]) );
  DFF_X1 \CWSE_reg[14]  ( .D(CWSD[14]), .CK(notClk), .Q(StatusMux81_sel[2]) );
  DFF_X1 \CWSF_reg2[16]  ( .D(n289), .CK(Clk), .Q(CWSF[16]) );
  DFF_X1 \CWSD_reg[16]  ( .D(CWSF[16]), .CK(notClk), .Q(CWSD[16]) );
  DFF_X1 \CWSE_reg[16]  ( .D(CWSD[16]), .CK(notClk), .Q(ALU_Unsign) );
  DFF_X1 \CWSF_reg2[18]  ( .D(n285), .CK(Clk), .Q(CWSF[18]) );
  DFF_X1 \CWSD_reg[18]  ( .D(CWSF[18]), .CK(notClk), .Q(CWSD[18]) );
  DFF_X1 \CWSE_reg[18]  ( .D(CWSD[18]), .CK(notClk), .Q(ALU_Sel[1]) );
  DFF_X1 \CWSF_reg2[20]  ( .D(n281), .CK(Clk), .Q(CWSF[20]) );
  DFF_X1 \CWSD_reg[20]  ( .D(CWSF[20]), .CK(notClk), .Q(CWSD[20]) );
  DFF_X1 \CWSE_reg[20]  ( .D(CWSD[20]), .CK(notClk), .Q(ALU_Sel[3]) );
  DFF_X1 \CWSF_reg2[22]  ( .D(n277), .CK(Clk), .Q(CWSF[22]) );
  DFF_X1 \CWSD_reg[22]  ( .D(CWSF[22]), .CK(notClk), .Q(CWSD[22]) );
  DFF_X1 \CWSF_reg2[24]  ( .D(n273), .CK(Clk), .Q(CWSF[24]) );
  DFF_X1 \CWSD_reg[24]  ( .D(CWSF[24]), .CK(notClk), .Q(CWSD[24]) );
  DFF_X1 \CWSF_reg2[26]  ( .D(n269), .CK(Clk), .Q(CWSF[26]) );
  DFF_X1 \CWSD_reg[26]  ( .D(CWSF[26]), .CK(notClk), .Q(ImmMux21_Sel) );
  DFF_X1 \CWSF_reg2[28]  ( .D(n266), .CK(Clk), .Q(CWSF[28]) );
  DFF_X1 \CWSD_reg[28]  ( .D(CWSF[28]), .CK(notClk), .Q(RWMux41WR_Sel[1]) );
  DFF_X1 \CWSF_reg2[30]  ( .D(n263), .CK(Clk), .Q(CWSF[30]) );
  DFF_X1 \CWSD_reg[30]  ( .D(CWSF[30]), .CK(notClk), .Q(R1Mux21A_Sel) );
  DFF_X1 \CWSF_reg2[32]  ( .D(n260), .CK(Clk), .Q(CWSF[32]) );
  DFF_X1 \CWSD_reg[32]  ( .D(CWSF[32]), .CK(notClk), .Q(RF_RD1) );
  DFF_X1 \CWSF_reg2[34]  ( .D(n257), .CK(Clk), .Q(CWSF[34]) );
  DFF_X1 \CWSF_reg2[36]  ( .D(n254), .CK(Clk), .Q(IRAM_Rst) );
  DFF_X1 \CWSF_reg2[38]  ( .D(n252), .CK(Clk), .Q(PCMux41_Sel[1]) );
  DFF_X1 \CWSF_reg2[40]  ( .D(n250), .CK(Clk), .Q(n784) );
  DFF_X1 JumpR_In_reg ( .D(n248), .CK(Clk), .Q(n753), .QN(n283) );
  DFF_X1 JumpRInst_reg ( .D(N3794), .CK(Clk), .Q(JumpRInst) );
  DFF_X1 LHIInst_reg ( .D(n246), .CK(Clk), .Q(LHIInst), .QN(n202) );
  DFF_X1 BranchZ_In_reg ( .D(n245), .CK(Clk), .Q(n711), .QN(n752) );
  DFF_X1 \CW_reg[38]  ( .D(n244), .CK(Clk), .Q(CW[38]) );
  DFF_X1 \CWSF_reg[38]  ( .D(CW[38]), .CK(notClk), .Q(PCMux41_Sel[1]) );
  DFF_X1 \CW_reg[37]  ( .D(n242), .CK(Clk), .Q(CW[37]) );
  DFF_X1 \CWSF_reg[37]  ( .D(CW[37]), .CK(notClk), .Q(PCMux41_Sel[0]) );
  DFF_X1 BranchInst_reg ( .D(n240), .CK(Clk), .Q(BranchInst), .QN(n199) );
  DFF_X1 \CWSD_reg[34]  ( .D(CWSF[34]), .CK(notClk), .Q(n785) );
  DFF_X1 \CWSD_reg[35]  ( .D(CWSF[35]), .CK(notClk), .Q(n786) );
  DFF_X1 \CWSF_reg[40]  ( .D(1'b1), .CK(notClk), .Q(n784) );
  DFF_X1 \CWSE_reg[25]  ( .D(CWSD[25]), .CK(notClk), .Q(n788) );
  DFF_X1 \CWSM_reg[11]  ( .D(CWSE[11]), .CK(notClk), .Q(n790) );
  DFF_X1 \CWSE_reg[24]  ( .D(CWSD[24]), .CK(notClk), .Q(n787) );
  DFF_X1 \CWSM_reg[10]  ( .D(CWSE[10]), .CK(notClk), .Q(n789) );
  DFF_X1 \CWSWB_reg[0]  ( .D(CWSM[0]), .CK(notClk), .Q(n792) );
  DFF_X2 \CWSE_reg[23]  ( .D(CWSD[23]), .CK(notClk), .Q(OPBMux41_Sel[1]) );
  DFF_X2 \CWSE_reg2[23]  ( .D(n489), .CK(Clk), .Q(OPBMux41_Sel[1]) );
  DFF_X1 Jump_reg ( .D(N3792), .CK(Clk), .Q(Jump) );
  INV_X2 U3 ( .A(Clk), .ZN(notClk) );
  NOR4_X2 U285 ( .A1(n251), .A2(n264), .A3(Inst[2]), .A4(Inst[3]), .ZN(n96) );
  NAND3_X1 U323 ( .A1(n57), .A2(n58), .A3(n59), .ZN(n628) );
  NAND3_X1 U324 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n65) );
  NAND3_X1 U325 ( .A1(n74), .A2(n75), .A3(n66), .ZN(n62) );
  NAND3_X1 U326 ( .A1(n84), .A2(Inst_28), .A3(n90), .ZN(n89) );
  NAND3_X1 U327 ( .A1(n84), .A2(n85), .A3(n101), .ZN(n100) );
  NAND3_X1 U328 ( .A1(n138), .A2(n120), .A3(n82), .ZN(n137) );
  NAND3_X1 U329 ( .A1(n164), .A2(n165), .A3(n771), .ZN(n163) );
  NAND3_X1 U330 ( .A1(n64), .A2(n164), .A3(n68), .ZN(n171) );
  NAND3_X1 U331 ( .A1(n66), .A2(n174), .A3(n68), .ZN(n172) );
  NAND3_X1 U332 ( .A1(n164), .A2(n105), .A3(n64), .ZN(n69) );
  NAND3_X1 U333 ( .A1(n93), .A2(n144), .A3(n152), .ZN(n179) );
  NAND3_X1 U334 ( .A1(n75), .A2(n185), .A3(n103), .ZN(n164) );
  NAND3_X1 U335 ( .A1(Inst_30), .A2(n198), .A3(n139), .ZN(n67) );
  NAND3_X1 U336 ( .A1(Inst_27), .A2(n75), .A3(n215), .ZN(n106) );
  NAND3_X1 U337 ( .A1(n198), .A2(n92), .A3(n243), .ZN(n105) );
  NAND3_X1 U338 ( .A1(n122), .A2(n253), .A3(n255), .ZN(n80) );
  NAND3_X1 U339 ( .A1(n152), .A2(n110), .A3(n261), .ZN(n123) );
  NAND3_X1 U340 ( .A1(n262), .A2(n256), .A3(n161), .ZN(n144) );
  NAND3_X1 U341 ( .A1(n259), .A2(Inst[5]), .A3(n148), .ZN(n265) );
  NAND3_X1 U342 ( .A1(n267), .A2(Inst[2]), .A3(n259), .ZN(n146) );
  NAND3_X1 U343 ( .A1(Inst[2]), .A2(n121), .A3(n267), .ZN(n147) );
  NAND3_X1 U344 ( .A1(n139), .A2(Inst_27), .A3(n215), .ZN(n70) );
  NAND3_X1 U345 ( .A1(Inst_28), .A2(n74), .A3(Inst_30), .ZN(n192) );
  NAND3_X1 U346 ( .A1(n198), .A2(n168), .A3(Inst_28), .ZN(n165) );
  NAND3_X1 U347 ( .A1(n243), .A2(n74), .A3(Inst_27), .ZN(n184) );
  DFF_X1 \CWSE_reg2[22]  ( .D(n487), .CK(Clk), .Q(OPBMux41_Sel[0]) );
  DFF_X1 \CWSE_reg[22]  ( .D(CWSD[22]), .CK(notClk), .Q(OPBMux41_Sel[0]) );
  DFF_X1 \CWSE_reg[21]  ( .D(CWSD[21]), .CK(notClk), .Q(OPAMux21_Sel) );
  DFF_X1 \CWSE_reg2[21]  ( .D(n485), .CK(Clk), .Q(OPAMux21_Sel) );
  NOR4_X1 U4 ( .A1(n168), .A2(n185), .A3(n170), .A4(Inst_28), .ZN(n134) );
  AND4_X1 U5 ( .A1(n192), .A2(n70), .A3(n193), .A4(n194), .ZN(n751) );
  INV_X1 U6 ( .A(n784), .ZN(n754) );
  INV_X16 U7 ( .A(n754), .ZN(FATCH_En) );
  CLKBUF_X3 U8 ( .A(n791), .Z(WBMux41_Sel[1]) );
  CLKBUF_X3 U9 ( .A(n789), .Z(MEMORY_Rst) );
  CLKBUF_X3 U10 ( .A(n787), .Z(EXECUTE_Rst) );
  INV_X1 U11 ( .A(n792), .ZN(n759) );
  INV_X8 U12 ( .A(n759), .ZN(WBMux41_Sel[0]) );
  INV_X1 U13 ( .A(n788), .ZN(n761) );
  INV_X8 U14 ( .A(n761), .ZN(EXECUTE_En) );
  INV_X1 U15 ( .A(n790), .ZN(n763) );
  INV_X8 U16 ( .A(n763), .ZN(MEMORY_En) );
  INV_X1 U17 ( .A(n785), .ZN(n765) );
  INV_X8 U18 ( .A(n765), .ZN(DECODE_Rst) );
  INV_X1 U19 ( .A(n786), .ZN(n767) );
  INV_X16 U20 ( .A(n767), .ZN(DECODE_En) );
  INV_X1 U21 ( .A(n69), .ZN(n66) );
  INV_X1 U22 ( .A(n58), .ZN(N3793) );
  INV_X1 U23 ( .A(n85), .ZN(n196) );
  NOR2_X1 U24 ( .A1(n53), .A2(n105), .ZN(n61) );
  INV_X1 U25 ( .A(n64), .ZN(n53) );
  INV_X1 U26 ( .A(n779), .ZN(n777) );
  NAND2_X1 U27 ( .A1(n63), .A2(n64), .ZN(n57) );
  INV_X1 U28 ( .A(n117), .ZN(n50) );
  AND3_X1 U29 ( .A1(n87), .A2(n777), .A3(n159), .ZN(n193) );
  INV_X1 U30 ( .A(n779), .ZN(n776) );
  INV_X1 U31 ( .A(n779), .ZN(n775) );
  INV_X1 U32 ( .A(n779), .ZN(n774) );
  NAND2_X1 U33 ( .A1(n109), .A2(n776), .ZN(n58) );
  NOR3_X1 U34 ( .A1(n63), .A2(n56), .A3(n197), .ZN(n85) );
  OAI21_X1 U35 ( .B1(n87), .B2(n139), .A(n52), .ZN(n197) );
  NAND2_X1 U36 ( .A1(n102), .A2(n139), .ZN(n159) );
  INV_X1 U37 ( .A(n144), .ZN(n132) );
  INV_X1 U38 ( .A(n115), .ZN(n120) );
  INV_X1 U39 ( .A(n158), .ZN(n149) );
  INV_X1 U40 ( .A(n78), .ZN(n162) );
  INV_X1 U41 ( .A(n113), .ZN(n262) );
  NOR2_X1 U42 ( .A1(n778), .A2(n751), .ZN(n64) );
  NAND4_X1 U43 ( .A1(n164), .A2(n105), .A3(n184), .A4(n774), .ZN(n117) );
  NAND2_X1 U44 ( .A1(n770), .A2(n166), .ZN(n180) );
  BUF_X1 U45 ( .A(n772), .Z(n779) );
  BUF_X1 U46 ( .A(n772), .Z(n780) );
  AND2_X1 U47 ( .A1(n777), .A2(n163), .ZN(n55) );
  BUF_X1 U48 ( .A(n772), .Z(n778) );
  OAI21_X1 U49 ( .B1(n774), .B2(n752), .A(n183), .ZN(n245) );
  NAND4_X1 U50 ( .A1(n49), .A2(n50), .A3(n92), .A4(n752), .ZN(n183) );
  AND4_X1 U51 ( .A1(n70), .A2(n105), .A3(n106), .A4(n107), .ZN(n84) );
  NOR3_X1 U52 ( .A1(n53), .A2(n108), .A3(n109), .ZN(n107) );
  NOR2_X1 U53 ( .A1(n184), .A2(n778), .ZN(N3792) );
  BUF_X1 U54 ( .A(n773), .Z(n783) );
  BUF_X1 U55 ( .A(n773), .Z(n782) );
  BUF_X1 U56 ( .A(n773), .Z(n781) );
  INV_X1 U57 ( .A(n181), .ZN(N3794) );
  AOI211_X1 U58 ( .C1(n162), .C2(n259), .A(n97), .B(n133), .ZN(n152) );
  AOI211_X1 U59 ( .C1(n121), .C2(n96), .A(n132), .B(n133), .ZN(n83) );
  NOR3_X1 U60 ( .A1(n168), .A2(n185), .A3(n275), .ZN(n102) );
  NOR4_X1 U61 ( .A1(n95), .A2(n96), .A3(n97), .A4(n98), .ZN(n94) );
  NOR2_X1 U62 ( .A1(n92), .A2(n75), .ZN(n139) );
  NOR3_X1 U63 ( .A1(n264), .A2(n258), .A3(n251), .ZN(n267) );
  AOI211_X1 U64 ( .C1(n96), .C2(n262), .A(n132), .B(n95), .ZN(n261) );
  AOI21_X1 U65 ( .B1(n75), .B2(n104), .A(n49), .ZN(n52) );
  NOR3_X1 U66 ( .A1(n112), .A2(n96), .A3(n97), .ZN(n111) );
  AOI21_X1 U67 ( .B1(n113), .B2(n114), .A(n115), .ZN(n112) );
  INV_X1 U68 ( .A(n96), .ZN(n79) );
  NAND2_X1 U69 ( .A1(n215), .A2(n170), .ZN(n87) );
  INV_X1 U70 ( .A(n165), .ZN(n49) );
  NOR2_X1 U71 ( .A1(n122), .A2(n138), .ZN(n113) );
  NOR2_X1 U72 ( .A1(n126), .A2(n185), .ZN(n158) );
  NAND2_X1 U73 ( .A1(n267), .A2(n256), .ZN(n78) );
  NAND4_X1 U74 ( .A1(n174), .A2(n200), .A3(n86), .A4(n106), .ZN(n124) );
  NAND2_X1 U75 ( .A1(n102), .A2(n103), .ZN(n200) );
  OAI21_X1 U76 ( .B1(n79), .B2(n131), .A(n83), .ZN(n129) );
  NAND2_X1 U77 ( .A1(n148), .A2(n264), .ZN(n115) );
  INV_X1 U78 ( .A(n70), .ZN(n73) );
  INV_X1 U79 ( .A(n253), .ZN(n251) );
  NAND2_X1 U80 ( .A1(n166), .A2(n175), .ZN(n109) );
  NAND2_X1 U81 ( .A1(n215), .A2(n103), .ZN(n86) );
  OAI21_X1 U82 ( .B1(n161), .B2(n162), .A(n138), .ZN(n160) );
  INV_X1 U83 ( .A(n134), .ZN(n140) );
  INV_X1 U84 ( .A(n67), .ZN(n63) );
  INV_X1 U85 ( .A(n147), .ZN(n97) );
  AND2_X1 U86 ( .A1(n146), .A2(n78), .ZN(n93) );
  INV_X1 U87 ( .A(n131), .ZN(n138) );
  INV_X1 U88 ( .A(n184), .ZN(n56) );
  INV_X1 U89 ( .A(n114), .ZN(n121) );
  INV_X1 U90 ( .A(n80), .ZN(n98) );
  INV_X1 U91 ( .A(n103), .ZN(n279) );
  AND2_X1 U92 ( .A1(n120), .A2(n259), .ZN(n95) );
  INV_X1 U93 ( .A(n91), .ZN(n126) );
  INV_X1 U94 ( .A(n108), .ZN(n174) );
  AND2_X1 U95 ( .A1(n175), .A2(n165), .ZN(n68) );
  AND2_X1 U96 ( .A1(n74), .A2(n170), .ZN(n198) );
  OR2_X1 U97 ( .A1(DECODE_En), .A2(n780), .ZN(n565) );
  OR2_X1 U98 ( .A1(n784), .A2(n780), .ZN(n250) );
  OR2_X1 U99 ( .A1(DECODE_Rst), .A2(n780), .ZN(n563) );
  OR2_X1 U100 ( .A1(MEMORY_En), .A2(n782), .ZN(n441) );
  OR2_X1 U101 ( .A1(EXECUTE_En), .A2(n781), .ZN(n493) );
  AND2_X1 U102 ( .A1(n777), .A2(WBMux41_Sel[0]), .ZN(n413) );
  OR2_X1 U103 ( .A1(EXECUTE_Rst), .A2(n781), .ZN(n491) );
  OR2_X1 U104 ( .A1(MEMORY_Rst), .A2(n782), .ZN(n439) );
  AND2_X1 U105 ( .A1(n777), .A2(WBMux41_Sel[1]), .ZN(n415) );
  AND2_X1 U106 ( .A1(OPBMux41_Sel[1]), .A2(n776), .ZN(n489) );
  AND2_X1 U107 ( .A1(RWMux41WR_Sel[0]), .A2(n774), .ZN(n549) );
  AND2_X1 U108 ( .A1(RWMux41WR_Sel[1]), .A2(n774), .ZN(n551) );
  AND2_X1 U109 ( .A1(R2Mux21B_Sel), .A2(n774), .ZN(n553) );
  AND2_X1 U110 ( .A1(R1Mux21A_Sel), .A2(n774), .ZN(n555) );
  OR2_X1 U111 ( .A1(CWSD[24]), .A2(n780), .ZN(n543) );
  OR2_X1 U112 ( .A1(RF_Rst), .A2(n780), .ZN(n561) );
  OR2_X1 U113 ( .A1(CWSF[34]), .A2(n783), .ZN(n257) );
  OR2_X1 U114 ( .A1(CWSF[24]), .A2(n783), .ZN(n273) );
  OR2_X1 U115 ( .A1(CWSF[10]), .A2(n783), .ZN(n302) );
  OR2_X1 U116 ( .A1(CWSF[8]), .A2(n783), .ZN(n307) );
  OR2_X1 U117 ( .A1(CWSF[11]), .A2(n783), .ZN(n360) );
  OR2_X1 U118 ( .A1(CWSF[25]), .A2(n783), .ZN(n388) );
  OR2_X1 U119 ( .A1(CWSF[33]), .A2(n783), .ZN(n400) );
  OR2_X1 U120 ( .A1(CWSF[35]), .A2(n782), .ZN(n403) );
  OR2_X1 U121 ( .A1(FS_Rst), .A2(n782), .ZN(n409) );
  OR2_X1 U122 ( .A1(DATAMEM_Rst), .A2(n782), .ZN(n435) );
  OR2_X1 U123 ( .A1(CWSE[8]), .A2(n782), .ZN(n459) );
  OR2_X1 U124 ( .A1(CWSE[10]), .A2(n781), .ZN(n463) );
  OR2_X1 U125 ( .A1(CWSE[11]), .A2(n781), .ZN(n465) );
  OR2_X1 U126 ( .A1(CWSD[8]), .A2(n782), .ZN(n511) );
  OR2_X1 U127 ( .A1(CWSD[10]), .A2(n781), .ZN(n515) );
  OR2_X1 U128 ( .A1(CWSD[11]), .A2(n781), .ZN(n517) );
  OR2_X1 U129 ( .A1(CWSD[25]), .A2(n781), .ZN(n545) );
  AND2_X1 U130 ( .A1(CWSF[12]), .A2(n776), .ZN(n297) );
  AND2_X1 U131 ( .A1(CWSF[6]), .A2(n776), .ZN(n312) );
  AND2_X1 U132 ( .A1(CWSF[4]), .A2(n776), .ZN(n317) );
  AND2_X1 U133 ( .A1(CWSF[2]), .A2(n776), .ZN(n323) );
  AND2_X1 U134 ( .A1(CWSF[0]), .A2(n776), .ZN(n329) );
  AND2_X1 U135 ( .A1(CWSF[1]), .A2(n776), .ZN(n335) );
  AND2_X1 U136 ( .A1(CWSF[3]), .A2(n776), .ZN(n340) );
  AND2_X1 U137 ( .A1(CWSF[5]), .A2(n776), .ZN(n345) );
  AND2_X1 U138 ( .A1(CWSF[7]), .A2(n776), .ZN(n350) );
  AND2_X1 U139 ( .A1(CWSF[9]), .A2(n776), .ZN(n355) );
  AND2_X1 U140 ( .A1(CWSF[13]), .A2(n776), .ZN(n364) );
  AND2_X1 U141 ( .A1(CWSF[15]), .A2(n776), .ZN(n368) );
  AND2_X1 U142 ( .A1(CWSF[17]), .A2(n776), .ZN(n372) );
  AND2_X1 U143 ( .A1(CWSF[19]), .A2(n776), .ZN(n376) );
  AND2_X1 U144 ( .A1(CWSF[21]), .A2(n776), .ZN(n380) );
  AND2_X1 U145 ( .A1(CWSF[23]), .A2(n776), .ZN(n384) );
  AND2_X1 U146 ( .A1(CWSF[27]), .A2(n776), .ZN(n391) );
  AND2_X1 U147 ( .A1(CWSF[29]), .A2(n776), .ZN(n394) );
  AND2_X1 U148 ( .A1(CWSF[31]), .A2(n776), .ZN(n397) );
  AND2_X1 U149 ( .A1(PCMux41_Sel[0]), .A2(n776), .ZN(n405) );
  AND2_X1 U150 ( .A1(FATCHRstMux21_Sel), .A2(n776), .ZN(n407) );
  AND2_X1 U151 ( .A1(RF_WR), .A2(n775), .ZN(n417) );
  AND2_X1 U152 ( .A1(CWSM[0]), .A2(n775), .ZN(n419) );
  AND2_X1 U153 ( .A1(CWSM[1]), .A2(n775), .ZN(n421) );
  AND2_X1 U154 ( .A1(CWSM[2]), .A2(n775), .ZN(n423) );
  AND2_X1 U155 ( .A1(DATAMEM_Unsign), .A2(n775), .ZN(n425) );
  AND2_X1 U156 ( .A1(DATAMEM_Byte), .A2(n775), .ZN(n427) );
  AND2_X1 U157 ( .A1(DATAMEM_HalfWord), .A2(n775), .ZN(n429) );
  AND2_X1 U158 ( .A1(DATAMEM_Word), .A2(n775), .ZN(n431) );
  AND2_X1 U159 ( .A1(DATAMEM_Read_Wrn), .A2(n775), .ZN(n433) );
  AND2_X1 U160 ( .A1(DATAMEM_En), .A2(n775), .ZN(n437) );
  AND2_X1 U161 ( .A1(CWSE[0]), .A2(n775), .ZN(n443) );
  AND2_X1 U162 ( .A1(CWSE[1]), .A2(n775), .ZN(n445) );
  AND2_X1 U163 ( .A1(CWSE[2]), .A2(n775), .ZN(n447) );
  AND2_X1 U164 ( .A1(CWSE[3]), .A2(n775), .ZN(n449) );
  AND2_X1 U165 ( .A1(CWSE[4]), .A2(n775), .ZN(n451) );
  AND2_X1 U166 ( .A1(CWSE[5]), .A2(n775), .ZN(n453) );
  AND2_X1 U167 ( .A1(CWSE[6]), .A2(n775), .ZN(n455) );
  AND2_X1 U168 ( .A1(CWSE[7]), .A2(n775), .ZN(n457) );
  AND2_X1 U169 ( .A1(CWSE[9]), .A2(n775), .ZN(n461) );
  AND2_X1 U170 ( .A1(StatusMux81_sel[0]), .A2(n775), .ZN(n467) );
  AND2_X1 U171 ( .A1(CWSD[13]), .A2(n775), .ZN(n521) );
  AND2_X1 U172 ( .A1(StatusMux81_sel[1]), .A2(n775), .ZN(n469) );
  AND2_X1 U173 ( .A1(StatusMux81_sel[2]), .A2(n776), .ZN(n471) );
  AND2_X1 U174 ( .A1(ALU_Arith_logN), .A2(n774), .ZN(n473) );
  AND2_X1 U175 ( .A1(ALU_Unsign), .A2(n775), .ZN(n475) );
  AND2_X1 U176 ( .A1(ALU_Sel[0]), .A2(n776), .ZN(n477) );
  AND2_X1 U177 ( .A1(ALU_Sel[1]), .A2(n775), .ZN(n479) );
  AND2_X1 U178 ( .A1(ALU_Sel[2]), .A2(n776), .ZN(n481) );
  AND2_X1 U179 ( .A1(ALU_Sel[3]), .A2(n775), .ZN(n483) );
  AND2_X1 U180 ( .A1(CWSD[0]), .A2(n776), .ZN(n495) );
  AND2_X1 U181 ( .A1(CWSD[1]), .A2(n775), .ZN(n497) );
  AND2_X1 U182 ( .A1(CWSD[2]), .A2(n776), .ZN(n499) );
  AND2_X1 U183 ( .A1(CWSD[3]), .A2(n775), .ZN(n501) );
  AND2_X1 U184 ( .A1(CWSD[4]), .A2(n776), .ZN(n503) );
  AND2_X1 U185 ( .A1(CWSD[5]), .A2(n775), .ZN(n505) );
  AND2_X1 U186 ( .A1(CWSD[6]), .A2(n776), .ZN(n507) );
  AND2_X1 U187 ( .A1(CWSD[7]), .A2(n775), .ZN(n509) );
  AND2_X1 U188 ( .A1(CWSD[9]), .A2(n776), .ZN(n513) );
  AND2_X1 U189 ( .A1(CWSD[12]), .A2(n775), .ZN(n519) );
  AND2_X1 U190 ( .A1(OPAMux21_Sel), .A2(n774), .ZN(n485) );
  AND2_X1 U191 ( .A1(PCMux41_Sel[1]), .A2(n777), .ZN(n252) );
  AND2_X1 U192 ( .A1(IRAM_Rst), .A2(n777), .ZN(n254) );
  AND2_X1 U193 ( .A1(CWSF[32]), .A2(n777), .ZN(n260) );
  AND2_X1 U194 ( .A1(CWSF[30]), .A2(n777), .ZN(n263) );
  AND2_X1 U195 ( .A1(CWSF[28]), .A2(n777), .ZN(n266) );
  AND2_X1 U196 ( .A1(CWSF[26]), .A2(n777), .ZN(n269) );
  AND2_X1 U197 ( .A1(CWSF[22]), .A2(n777), .ZN(n277) );
  AND2_X1 U198 ( .A1(CWSF[20]), .A2(n777), .ZN(n281) );
  AND2_X1 U199 ( .A1(CWSF[18]), .A2(n777), .ZN(n285) );
  AND2_X1 U200 ( .A1(CWSF[16]), .A2(n777), .ZN(n289) );
  AND2_X1 U201 ( .A1(CWSF[14]), .A2(n777), .ZN(n293) );
  AND2_X1 U202 ( .A1(CWSD[14]), .A2(n774), .ZN(n523) );
  AND2_X1 U203 ( .A1(CWSD[15]), .A2(n774), .ZN(n525) );
  AND2_X1 U204 ( .A1(CWSD[16]), .A2(n774), .ZN(n527) );
  AND2_X1 U205 ( .A1(CWSD[17]), .A2(n774), .ZN(n529) );
  AND2_X1 U206 ( .A1(CWSD[18]), .A2(n774), .ZN(n531) );
  AND2_X1 U207 ( .A1(CWSD[19]), .A2(n774), .ZN(n533) );
  AND2_X1 U208 ( .A1(CWSD[20]), .A2(n774), .ZN(n535) );
  AND2_X1 U209 ( .A1(CWSD[21]), .A2(n774), .ZN(n537) );
  AND2_X1 U210 ( .A1(CWSD[22]), .A2(n774), .ZN(n539) );
  AND2_X1 U211 ( .A1(CWSD[23]), .A2(n774), .ZN(n541) );
  AND2_X1 U212 ( .A1(ImmMux21_Sel), .A2(n774), .ZN(n547) );
  AND2_X1 U213 ( .A1(RF_RD2), .A2(n774), .ZN(n557) );
  AND2_X1 U214 ( .A1(RF_RD1), .A2(n774), .ZN(n559) );
  NOR3_X1 U215 ( .A1(n159), .A2(Inst_27), .A3(n53), .ZN(n130) );
  OAI222_X1 U216 ( .A1(n116), .A2(n117), .B1(n118), .B2(n119), .C1(n220), .C2(
        n770), .ZN(n601) );
  NOR3_X1 U217 ( .A1(n124), .A2(n63), .A3(n125), .ZN(n116) );
  AOI221_X1 U218 ( .B1(n120), .B2(n121), .C1(n122), .C2(Inst[5]), .A(n123), 
        .ZN(n118) );
  INV_X1 U219 ( .A(n61), .ZN(n119) );
  NOR3_X1 U220 ( .A1(n53), .A2(Inst_28), .A3(n149), .ZN(n143) );
  OAI221_X1 U221 ( .B1(n69), .B2(n70), .C1(n226), .C2(n771), .A(n62), .ZN(n613) );
  NAND4_X1 U222 ( .A1(n64), .A2(Inst_31), .A3(n170), .A4(n168), .ZN(n169) );
  OAI221_X1 U223 ( .B1(n53), .B2(n149), .C1(n216), .C2(n771), .A(n150), .ZN(
        n593) );
  AOI21_X1 U224 ( .B1(n61), .B2(n151), .A(n130), .ZN(n150) );
  OAI211_X1 U225 ( .C1(n114), .C2(n78), .A(n146), .B(n152), .ZN(n151) );
  OAI221_X1 U226 ( .B1(n53), .B2(n140), .C1(n217), .C2(n770), .A(n141), .ZN(
        n595) );
  AOI21_X1 U227 ( .B1(n82), .B2(n142), .A(n143), .ZN(n141) );
  NAND2_X1 U228 ( .A1(n78), .A2(n144), .ZN(n142) );
  OAI221_X1 U229 ( .B1(n53), .B2(n136), .C1(n218), .C2(n770), .A(n137), .ZN(
        n597) );
  NAND2_X1 U230 ( .A1(n104), .A2(n139), .ZN(n136) );
  OAI221_X1 U231 ( .B1(n127), .B2(n53), .C1(n219), .C2(n771), .A(n128), .ZN(
        n599) );
  AOI221_X1 U232 ( .B1(n134), .B2(Inst_31), .C1(Inst_26), .C2(n135), .A(n73), 
        .ZN(n127) );
  AOI21_X1 U233 ( .B1(n82), .B2(n129), .A(n130), .ZN(n128) );
  OAI21_X1 U234 ( .B1(Inst_28), .B2(n87), .A(n106), .ZN(n135) );
  OAI221_X1 U235 ( .B1(n52), .B2(n53), .C1(n238), .C2(n771), .A(n54), .ZN(n639) );
  INV_X1 U236 ( .A(N3792), .ZN(n54) );
  OAI221_X1 U237 ( .B1(Inst_26), .B2(n153), .C1(n295), .C2(n770), .A(n154), 
        .ZN(n591) );
  INV_X1 U238 ( .A(n143), .ZN(n153) );
  AOI211_X1 U239 ( .C1(n61), .C2(n155), .A(n130), .B(n156), .ZN(n154) );
  NAND2_X1 U240 ( .A1(n152), .A2(n160), .ZN(n155) );
  NOR3_X1 U241 ( .A1(n53), .A2(n157), .A3(n92), .ZN(n156) );
  AOI21_X1 U242 ( .B1(n158), .B2(Inst_28), .A(n134), .ZN(n157) );
  OAI211_X1 U243 ( .C1(n204), .C2(n770), .A(n172), .B(n173), .ZN(n569) );
  NAND4_X1 U244 ( .A1(n61), .A2(n152), .A3(n93), .A4(n144), .ZN(n173) );
  OAI211_X1 U245 ( .C1(n221), .C2(n771), .A(n99), .B(n100), .ZN(n603) );
  NAND4_X1 U246 ( .A1(n61), .A2(n110), .A3(n83), .A4(n111), .ZN(n99) );
  AOI21_X1 U247 ( .B1(n102), .B2(n103), .A(n104), .ZN(n101) );
  OAI211_X1 U248 ( .C1(n222), .C2(n771), .A(n88), .B(n89), .ZN(n605) );
  NAND4_X1 U249 ( .A1(n61), .A2(n93), .A3(n83), .A4(n94), .ZN(n88) );
  AOI21_X1 U250 ( .B1(n91), .B2(n92), .A(n49), .ZN(n90) );
  OAI211_X1 U251 ( .C1(n230), .C2(n771), .A(n62), .B(n57), .ZN(n622) );
  OAI22_X1 U252 ( .A1(n210), .A2(n770), .B1(n53), .B2(n166), .ZN(n581) );
  OAI22_X1 U253 ( .A1(n206), .A2(n770), .B1(n75), .B2(n169), .ZN(n573) );
  OAI22_X1 U254 ( .A1(n207), .A2(n770), .B1(Inst_26), .B2(n169), .ZN(n575) );
  OAI22_X1 U255 ( .A1(n208), .A2(n770), .B1(n92), .B2(n169), .ZN(n577) );
  OAI22_X1 U256 ( .A1(n234), .A2(n770), .B1(n56), .B2(n53), .ZN(n630) );
  OAI22_X1 U257 ( .A1(n709), .A2(n778), .B1(n711), .B2(n191), .ZN(n242) );
  AOI221_X1 U258 ( .B1(n775), .B2(n753), .C1(n751), .C2(CW[37]), .A(N3792), 
        .ZN(n191) );
  OAI21_X1 U259 ( .B1(n228), .B2(n770), .A(n55), .ZN(n617) );
  OAI21_X1 U260 ( .B1(n229), .B2(n770), .A(n65), .ZN(n620) );
  OAI21_X1 U261 ( .B1(n232), .B2(n770), .A(n57), .ZN(n626) );
  OAI21_X1 U262 ( .B1(n235), .B2(n770), .A(n774), .ZN(n632) );
  OAI21_X1 U263 ( .B1(n236), .B2(n770), .A(n774), .ZN(n634) );
  OAI21_X1 U264 ( .B1(n237), .B2(n770), .A(n55), .ZN(n636) );
  OAI21_X1 U265 ( .B1(n239), .B2(n770), .A(n774), .ZN(n642) );
  OAI21_X1 U266 ( .B1(n205), .B2(n771), .A(n171), .ZN(n571) );
  OAI21_X1 U267 ( .B1(n209), .B2(n771), .A(n167), .ZN(n579) );
  NAND4_X1 U268 ( .A1(n64), .A2(Inst_31), .A3(Inst_27), .A4(n168), .ZN(n167)
         );
  OAI21_X1 U269 ( .B1(n211), .B2(n771), .A(n774), .ZN(n583) );
  OAI21_X1 U270 ( .B1(n212), .B2(n771), .A(n58), .ZN(n585) );
  OAI21_X1 U271 ( .B1(n213), .B2(n771), .A(n774), .ZN(n587) );
  OAI21_X1 U272 ( .B1(n214), .B2(n771), .A(n55), .ZN(n589) );
  OAI21_X1 U273 ( .B1(n224), .B2(n771), .A(n62), .ZN(n609) );
  OAI21_X1 U274 ( .B1(n225), .B2(n771), .A(n71), .ZN(n611) );
  NAND4_X1 U275 ( .A1(n50), .A2(n771), .A3(n72), .A4(n67), .ZN(n71) );
  NOR2_X1 U276 ( .A1(n49), .A2(n73), .ZN(n72) );
  OAI21_X1 U277 ( .B1(n227), .B2(n771), .A(n774), .ZN(n615) );
  OAI21_X1 U278 ( .B1(n231), .B2(n771), .A(n57), .ZN(n624) );
  NOR4_X1 U279 ( .A1(n195), .A2(n124), .A3(n109), .A4(n196), .ZN(n194) );
  OAI211_X1 U280 ( .C1(n223), .C2(n770), .A(n76), .B(n77), .ZN(n607) );
  NAND4_X1 U281 ( .A1(n84), .A2(n85), .A3(n86), .A4(n87), .ZN(n76) );
  NAND4_X1 U282 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .ZN(n77) );
  AND2_X1 U283 ( .A1(n82), .A2(n83), .ZN(n81) );
  AOI21_X1 U284 ( .B1(n53), .B2(n176), .A(n177), .ZN(n567) );
  NAND2_X1 U286 ( .A1(n774), .A2(CW[0]), .ZN(n176) );
  AOI211_X1 U287 ( .C1(n178), .C2(n179), .A(n180), .B(n108), .ZN(n177) );
  INV_X1 U288 ( .A(n105), .ZN(n178) );
  OAI21_X1 U289 ( .B1(n709), .B2(n775), .A(n48), .ZN(n643) );
  NAND4_X1 U290 ( .A1(n709), .A2(Inst_26), .A3(n49), .A4(n50), .ZN(n48) );
  AND4_X1 U291 ( .A1(n61), .A2(n145), .A3(n146), .A4(n147), .ZN(n82) );
  NAND2_X1 U292 ( .A1(n148), .A2(Inst[5]), .ZN(n145) );
  OAI21_X1 U293 ( .B1(n753), .B2(n187), .A(n188), .ZN(n244) );
  INV_X1 U294 ( .A(n189), .ZN(n188) );
  NAND2_X1 U295 ( .A1(n751), .A2(CW[38]), .ZN(n187) );
  AOI21_X1 U296 ( .B1(n752), .B2(n709), .A(n779), .ZN(n189) );
  AOI21_X1 U297 ( .B1(n751), .B2(CW[31]), .A(n61), .ZN(n59) );
  BUF_X1 U298 ( .A(Rst), .Z(n772) );
  OAI22_X1 U299 ( .A1(n202), .A2(n776), .B1(n779), .B2(n70), .ZN(n246) );
  NAND4_X1 U300 ( .A1(n283), .A2(n104), .A3(n75), .A4(n774), .ZN(n181) );
  OAI21_X1 U301 ( .B1(n199), .B2(n775), .A(n276), .ZN(n240) );
  OAI211_X1 U302 ( .C1(n278), .C2(N3794), .A(n752), .B(n709), .ZN(n276) );
  NOR3_X1 U303 ( .A1(n753), .A2(n778), .A3(n165), .ZN(n278) );
  OAI21_X1 U304 ( .B1(n283), .B2(n776), .A(n181), .ZN(n248) );
  BUF_X1 U305 ( .A(Rst), .Z(n773) );
  NOR3_X1 U306 ( .A1(n256), .A2(Inst[3]), .A3(n251), .ZN(n148) );
  NOR3_X1 U307 ( .A1(Inst_30), .A2(Inst_31), .A3(n185), .ZN(n215) );
  NOR4_X1 U308 ( .A1(Inst[4]), .A2(Inst[6]), .A3(Inst[10]), .A4(n274), .ZN(
        n253) );
  OR3_X1 U309 ( .A1(Inst[7]), .A2(Inst[9]), .A3(Inst[8]), .ZN(n274) );
  NOR2_X1 U310 ( .A1(n170), .A2(Inst_26), .ZN(n103) );
  NOR3_X1 U311 ( .A1(Inst_27), .A2(Inst_31), .A3(n168), .ZN(n91) );
  OAI211_X1 U312 ( .C1(Inst_27), .C2(n159), .A(n140), .B(n149), .ZN(n108) );
  NOR2_X1 U313 ( .A1(Inst[0]), .A2(Inst[1]), .ZN(n259) );
  AOI211_X1 U314 ( .C1(n87), .C2(n126), .A(n75), .B(Inst_26), .ZN(n125) );
  NOR2_X1 U315 ( .A1(n272), .A2(Inst[0]), .ZN(n122) );
  INV_X1 U316 ( .A(Inst_30), .ZN(n168) );
  NOR2_X1 U317 ( .A1(Inst_31), .A2(Inst_29), .ZN(n74) );
  INV_X1 U318 ( .A(Inst_28), .ZN(n75) );
  NAND4_X1 U319 ( .A1(n185), .A2(n168), .A3(n279), .A4(n282), .ZN(n166) );
  AOI21_X1 U320 ( .B1(Inst_27), .B2(Inst_28), .A(n275), .ZN(n282) );
  NOR3_X1 U321 ( .A1(n256), .A2(Inst[5]), .A3(n258), .ZN(n255) );
  INV_X1 U322 ( .A(Inst_26), .ZN(n92) );
  INV_X1 U348 ( .A(Inst_29), .ZN(n185) );
  NOR2_X1 U349 ( .A1(Inst_30), .A2(Inst_28), .ZN(n243) );
  AOI21_X1 U350 ( .B1(n233), .B2(n241), .A(n105), .ZN(n195) );
  AOI211_X1 U351 ( .C1(n138), .C2(n120), .A(n98), .B(n249), .ZN(n241) );
  AOI221_X1 U352 ( .B1(n96), .B2(n259), .C1(n122), .C2(n148), .A(n123), .ZN(
        n233) );
  NOR3_X1 U353 ( .A1(n251), .A2(Inst[3]), .A3(n114), .ZN(n249) );
  INV_X1 U354 ( .A(Inst_27), .ZN(n170) );
  NAND2_X1 U355 ( .A1(Inst[0]), .A2(n272), .ZN(n114) );
  AND3_X1 U356 ( .A1(Inst_27), .A2(n74), .A3(Inst_30), .ZN(n104) );
  NAND4_X1 U357 ( .A1(Inst_31), .A2(Inst_29), .A3(n243), .A4(n279), .ZN(n175)
         );
  INV_X1 U358 ( .A(Inst[5]), .ZN(n264) );
  INV_X1 U359 ( .A(Inst[2]), .ZN(n256) );
  INV_X1 U360 ( .A(Inst[3]), .ZN(n258) );
  AND3_X1 U361 ( .A1(n121), .A2(n161), .A3(Inst[2]), .ZN(n133) );
  NAND2_X1 U362 ( .A1(Inst[1]), .A2(Inst[0]), .ZN(n131) );
  AND2_X1 U363 ( .A1(n268), .A2(n270), .ZN(n161) );
  NOR4_X1 U364 ( .A1(Inst[10]), .A2(n258), .A3(n271), .A4(n264), .ZN(n268) );
  NOR4_X1 U365 ( .A1(Inst[9]), .A2(Inst[8]), .A3(Inst[7]), .A4(Inst[6]), .ZN(
        n270) );
  INV_X1 U366 ( .A(Inst[4]), .ZN(n271) );
  INV_X1 U370 ( .A(Inst[1]), .ZN(n272) );
  INV_X1 U371 ( .A(Inst_31), .ZN(n275) );
  AND2_X1 U372 ( .A1(n93), .A2(n265), .ZN(n110) );
  CLKBUF_X1 U373 ( .A(OPBMux41_Sel[0]), .Z(n769) );
  AND2_X1 U374 ( .A1(n769), .A2(n776), .ZN(n487) );
  INV_X1 U375 ( .A(n751), .ZN(n770) );
  INV_X1 U376 ( .A(n751), .ZN(n771) );
endmodule



    module datapath_Nbit32_RAM_DEPTH30_I_SIZE32_DATA_MEM_SIZE10_Nlogicfun3_NALUop4 ( 
        Rst, Clk, Inst, BrNZ, BrZ, BranchInst, StoreInst, JumpRInst, LHIInst, 
        FS_Rst, FATCHRstMux21_Sel, FATCH_En, PCMux41_Sel, Jump, IRAM_Rst, 
        DECODE_Rst, DECODE_En, RF_Rst, RF_RD1, RF_RD2, R1Mux21A_Sel, 
        R2Mux21B_Sel, RWMux41WR_Sel, ImmMux21_Sel, EXECUTE_Rst, EXECUTE_En, 
        OPAMux21_Sel, OPBMux41_Sel, ALU_Sel, ALU_Unsign, ALU_Arith_logN, 
        StatusMux81_sel, MEMORY_Rst, MEMORY_En, DATAMEM_En, DATAMEM_Rst, 
        DATAMEM_Read_Wrn, DATAMEM_Word, DATAMEM_HalfWord, DATAMEM_Byte, 
        DATAMEM_Unsign, RF_WR, WBMux41_Sel );
  output [31:0] Inst;
  input [1:0] PCMux41_Sel;
  input [1:0] RWMux41WR_Sel;
  input [1:0] OPBMux41_Sel;
  input [3:0] ALU_Sel;
  input [2:0] StatusMux81_sel;
  input [1:0] WBMux41_Sel;
  input Rst, Clk, BranchInst, StoreInst, JumpRInst, LHIInst, FS_Rst,
         FATCHRstMux21_Sel, FATCH_En, Jump, IRAM_Rst, DECODE_Rst, DECODE_En,
         RF_Rst, RF_RD1, RF_RD2, R1Mux21A_Sel, R2Mux21B_Sel, ImmMux21_Sel,
         EXECUTE_Rst, EXECUTE_En, OPAMux21_Sel, ALU_Unsign, ALU_Arith_logN,
         MEMORY_Rst, MEMORY_En, DATAMEM_En, DATAMEM_Rst, DATAMEM_Read_Wrn,
         DATAMEM_Word, DATAMEM_HalfWord, DATAMEM_Byte, DATAMEM_Unsign, RF_WR;
  output BrNZ, BrZ;
  wire   NPCReg_Rst, Branch_DO, JRInst_Del, FATCHRst_DO, StoreInstDel,
         \WB_Status[0] , Jump_DO, LHIInst_DEC, StoreInstEX, LHIInst_EXE,
         ALU_AeqB, ALU_AnoteqB, ALU_AgB, ALU_AlB, ALU_AgeqB, ALU_AleqB, Status,
         StoreInstMEM, StatusMEM, net291429;
  wire   [10:0] IRReg_Out;
  wire   [4:0] RF_AddrR1;
  wire   [4:0] RF_AddrR2;
  wire   [4:0] RF_AddrR3;
  wire   [25:0] ImmediateJ;
  wire   [31:26] IRReg_0_Out;
  wire   [31:16] ALU_opImm;
  wire   [31:16] LHI_Num;
  wire   [31:0] MEM_DataIn;
  wire   [4:0] RF_AddrWR;
  wire   [31:0] PC_Up;
  wire   [31:0] PC_Next;
  wire   [31:0] PC_New;
  wire   [31:0] PC_Datapath;
  wire   [29:0] PC_Inst;
  wire   [31:0] PC_Branch_Del;
  wire   [31:0] PC_Now;
  wire   [31:0] PC_Branch;
  wire   [31:0] PC_Actual;
  wire   [31:0] JumpAddr;
  wire   [29:0] IRAM_Addr;
  wire   [29:0] Addr_IRAM;
  wire   [31:0] NPCReg_Out;
  wire   [4:0] RF_AddrRD1;
  wire   [4:0] RF_AddrRD2;
  wire   [4:0] RF_AddrWRR3;
  wire   [31:0] RF_DataIn;
  wire   [31:0] ImmediateIop_ex;
  wire   [31:0] ImmediateI_ex;
  wire   [31:0] ImmediateJ_ex;
  wire   [31:0] Immediate;
  wire   [31:0] PC_BranchAdd;
  wire   [31:0] ALU_opA;
  wire   [31:0] ALU_opB;
  wire   [4:0] RF_WrAddr_EX;
  wire   [31:0] PC_Ret_Del;
  wire   [31:0] PC_Ret;
  wire   [31:0] ALU_Op1;
  wire   [31:0] Op2;
  wire   [31:0] Op1;
  wire   [31:0] ALU_Out;
  wire   [31:0] MEM_Addr;
  wire   [4:0] RF_WrAddr_MEM;
  wire   [31:0] Data_MEM_DataIn;
  wire   [9:0] Data_MEM_Addr;
  wire   [31:0] MEM_DataOut;
  wire   [31:0] WB_MEM;
  wire   [31:0] WB_ALU;
  tri   [1:0] PCMux41_Sel;
  tri   RF_RD1;
  tri   RF_RD2;
  tri   R1Mux21A_Sel;
  tri   R2Mux21B_Sel;
  tri   [1:0] RWMux41WR_Sel;
  tri   OPAMux21_Sel;
  tri   \OPBMux41_Sel[1] ;
  tri   [3:0] ALU_Sel;
  tri   ALU_Unsign;
  tri   ALU_Arith_logN;
  tri   [2:0] StatusMux81_sel;
  tri   DATAMEM_En;
  tri   DATAMEM_Rst;
  tri   DATAMEM_Read_Wrn;
  tri   DATAMEM_Word;
  tri   DATAMEM_HalfWord;
  tri   DATAMEM_Byte;
  tri   DATAMEM_Unsign;
  tri   RF_WR;
  tri   [31:0] RF_Out1;
  tri   [31:0] RF_Out2;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27;
  assign net291429 = OPBMux41_Sel[0];

  mux21N_N32_0 BrPCNextMux21 ( .in1(PC_Up), .in0(PC_Next), .S(Branch_DO), .U(
        PC_New) );
  PC_RAM_DEPTH30 PCinst ( .PC_In(PC_New), .En(FATCH_En), .Clk(Clk), .Res(Rst), 
        .PC_DATAP(PC_Datapath), .PC_IRAM(PC_Inst) );
  mux21N_N32_16 BrPCAddMux21 ( .in1(PC_Branch_Del), .in0(PC_Datapath), .S(
        Branch_DO), .U(PC_Now) );
  MUX21_40 JumpSel ( .in1(1'b1), .in0(Jump), .S(JRInst_Del), .Y(Jump_DO) );
  mux21N_N32_15 JmPCAddMux21 ( .in1(PC_Branch), .in0(PC_Now), .S(Jump_DO), .U(
        PC_Actual) );
  AddSubN_Nbit32_0 PCAdd ( .A(PC_Actual), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .addnsub(1'b0), .S(PC_Up) );
  FD_EN_0 jumpRFF ( .D(JumpRInst), .Clk(Clk), .RESET(1'b0), .EN(1'b1), .Q(
        JRInst_Del) );
  mux41 PCMux41sel ( .in3(BrNZ), .in2(BrZ), .in1(1'b0), .in0(1'b0), .sel(
        PCMux41_Sel), .Y(Branch_DO) );
  MUX21_800 FATCHRstMux21 ( .in1(1'b1), .in0(Rst), .S(FATCHRst_DO), .Y(
        NPCReg_Rst) );
  RegEn_Nbit32_0 BranchReg ( .A(PC_Branch), .Clk(Clk), .Reset(1'b0), .EN(1'b1), 
        .U(PC_Branch_Del) );
  mux21N_N32_14 BrAddrMux21 ( .in1(PC_Branch_Del), .in0(PC_Branch), .S(
        Branch_DO), .U(JumpAddr) );
  mux21N_N32_13 PCMux21 ( .in1(JumpAddr), .in0(PC_Up), .S(Branch_DO), .U(
        PC_Next) );
  mux21N_N30_0 AddrIRAMMux21 ( .in1(PC_Next[31:2]), .in0(PC_Inst), .S(
        Branch_DO), .U(IRAM_Addr) );
  mux21N_N30_1 JmAddrIRAMMux21 ( .in1(PC_Branch[31:2]), .in0(IRAM_Addr), .S(
        Jump_DO), .U(Addr_IRAM) );
  IRAM IRAMinst ( .Rst(Rst), .Addr(Addr_IRAM), .Dout(Inst) );
  FD_EN_438 StoreFF ( .D(StoreInst), .Clk(Clk), .RESET(NPCReg_Rst), .EN(1'b1), 
        .Q(StoreInstDel) );
  RegEn_Nbit32_12 NPCReg ( .A(PC_Next), .Clk(Clk), .Reset(1'b0), .EN(FATCH_En), 
        .U(NPCReg_Out) );
  RegEn_Nbit32_11 IRReg_0 ( .A(Inst), .Clk(Clk), .Reset(Rst), .EN(FATCH_En), 
        .U({IRReg_0_Out, ImmediateJ}) );
  RegEn_Nbit32_10 IRReg_1 ( .A({IRReg_0_Out, ImmediateJ}), .Clk(Clk), .Reset(
        NPCReg_Rst), .EN(FATCH_En), .U({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, RF_AddrR1, RF_AddrR2, RF_AddrR3, IRReg_Out})
         );
  FD_EN_437 LHIFFIF ( .D(LHIInst), .Clk(Clk), .RESET(NPCReg_Rst), .EN(1'b1), 
        .Q(LHIInst_DEC) );
  mux21N_N5_8 R1Mux21A ( .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in0(RF_AddrR1), 
        .S(R1Mux21A_Sel), .U(RF_AddrRD1) );
  mux21N_N5_36 R2Mux21B ( .in1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in0(RF_AddrR2), .S(R2Mux21B_Sel), .U(RF_AddrRD2) );
  mux41N_Nbit5 RWMux41WR ( .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in2({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .in1(RF_AddrR2), .in0(RF_AddrR3), .sel(
        RWMux41WR_Sel), .Y(RF_AddrWRR3) );
  register_file_Nbit32 RF ( .CLK(Clk), .RESET(Rst), .ENABLE(1'b1), .RD1(RF_RD1), .RD2(RF_RD2), .WR(RF_WR), .ADD_WR(RF_AddrWR), .ADD_RD1(RF_AddrRD1), 
        .ADD_RD2(RF_AddrRD2), .DATAIN(RF_DataIn), .OUT1(RF_Out1), .OUT2(
        RF_Out2) );
  signExtension_Nbitin16_Nbitout32_0 signex16I ( .A({RF_AddrR3, IRReg_Out}), 
        .Aextended(ImmediateIop_ex) );
  signExtension_Nbitin16_Nbitout32_1 signex16 ( .A(ImmediateJ[15:0]), 
        .Aextended(ImmediateI_ex) );
  signExtension_Nbitin26_Nbitout32 signex26 ( .A(ImmediateJ), .Aextended(
        ImmediateJ_ex) );
  AddSubN_Nbit32_2 BranchAdd ( .A(NPCReg_Out), .B(Immediate), .addnsub(1'b0), 
        .S(PC_BranchAdd) );
  mux21N_N32_12 JRMux21 ( .in1(RF_Out1), .in0(PC_BranchAdd), .S(JRInst_Del), 
        .U(PC_Branch) );
  zerotest_Nbit32 zero ( .A(RF_Out1), .zero(BrZ) );
  mux21N_N32_11 ImmMux21 ( .in1(ImmediateJ_ex), .in0(ImmediateI_ex), .S(Jump), 
        .U(Immediate) );
  FD_EN_436 StoreFFEX ( .D(StoreInstDel), .Clk(Clk), .RESET(DECODE_Rst), .EN(
        1'b1), .Q(StoreInstEX) );
  RegEn_Nbit32_9 AReg ( .A(RF_Out1), .Clk(Clk), .Reset(DECODE_Rst), .EN(
        DECODE_En), .U(ALU_opA) );
  RegEn_Nbit32_8 BReg ( .A(RF_Out2), .Clk(Clk), .Reset(DECODE_Rst), .EN(
        DECODE_En), .U(ALU_opB) );
  RegEn_Nbit32_7 ImmReg ( .A(ImmediateIop_ex), .Clk(Clk), .Reset(DECODE_Rst), 
        .EN(DECODE_En), .U({ALU_opImm, LHI_Num}) );
  RegEn_Nbit5_0 RFWRAddrID ( .A(RF_AddrWRR3), .Clk(Clk), .Reset(DECODE_Rst), 
        .EN(DECODE_En), .U(RF_WrAddr_EX) );
  RegEn_Nbit32_6 DelPCRetReg ( .A(NPCReg_Out), .Clk(Clk), .Reset(DECODE_Rst), 
        .EN(1'b1), .U(PC_Ret_Del) );
  RegEn_Nbit32_5 PCRetReg ( .A(PC_Ret_Del), .Clk(Clk), .Reset(DECODE_Rst), 
        .EN(DECODE_En), .U(PC_Ret) );
  FD_EN_435 LHIFFID ( .D(LHIInst_DEC), .Clk(Clk), .RESET(DECODE_Rst), .EN(1'b1), .Q(LHIInst_EXE) );
  mux21N_N32_10 OPAMux21 ( .in1(PC_Ret), .in0(ALU_opA), .S(OPAMux21_Sel), .U(
        ALU_Op1) );
  mux41N_Nbit32_0 OPBMux41 ( .in3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .in2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .in1({ALU_opImm, LHI_Num}), .in0(ALU_opB), .sel({OPBMux41_Sel[1], 
        net291429}), .Y(Op2) );
  mux21N_N32_9 OPALHIMux21 ( .in1({LHI_Num, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .in0(
        ALU_Op1), .S(LHIInst_EXE), .U(Op1) );
  ALU_v2 ALU ( .A(Op1), .B(Op2), .ALUsel(ALU_Sel), .unsign(ALU_Unsign), 
        .arith_logN(ALU_Arith_logN), .ALUout(ALU_Out), .AeqB(ALU_AeqB), 
        .AnoteqB(ALU_AnoteqB), .AgB(ALU_AgB), .AlB(ALU_AlB), .AgeqB(ALU_AgeqB), 
        .AleqB(ALU_AleqB) );
  mux81 StatusMux81 ( .in7(ALU_AeqB), .in6(ALU_AnoteqB), .in5(ALU_AgB), .in4(
        ALU_AlB), .in3(ALU_AgeqB), .in2(ALU_AleqB), .in1(1'b0), .in0(1'b0), 
        .sel(StatusMux81_sel), .Y(Status) );
  FD_EN_434 StoreFFMEM ( .D(StoreInstEX), .Clk(Clk), .RESET(EXECUTE_Rst), .EN(
        1'b1), .Q(StoreInstMEM) );
  RegEn_Nbit32_4 ALUReg ( .A(ALU_Out), .Clk(Clk), .Reset(EXECUTE_Rst), .EN(
        EXECUTE_En), .U(MEM_DataIn) );
  RegEn_Nbit32_3 DMEMAddrReg ( .A(ALU_opB), .Clk(Clk), .Reset(EXECUTE_Rst), 
        .EN(EXECUTE_En), .U(MEM_Addr) );
  RegEn_Nbit5_2 RFWRAddrEX ( .A(RF_WrAddr_EX), .Clk(Clk), .Reset(EXECUTE_Rst), 
        .EN(EXECUTE_En), .U(RF_WrAddr_MEM) );
  FD_EN_433 StatusRegEX ( .D(Status), .Clk(Clk), .RESET(EXECUTE_Rst), .EN(
        EXECUTE_En), .Q(StatusMEM) );
  mux21N_N32_8 SDATAMux21 ( .in1(MEM_Addr), .in0(MEM_DataIn), .S(StoreInstMEM), 
        .U(Data_MEM_DataIn) );
  mux21N_N32_7 SADDMux21 ( .in1(MEM_DataIn), .in0(MEM_Addr), .S(StoreInstMEM), 
        .U({SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, Data_MEM_Addr}) );
  DataMemory DataMem ( .DataIn(Data_MEM_DataIn), .Addr(Data_MEM_Addr), .En(
        DATAMEM_En), .Clk(Clk), .Rst(DATAMEM_Rst), .Read_Wrn(DATAMEM_Read_Wrn), 
        .Word(DATAMEM_Word), .HalfWord(DATAMEM_HalfWord), .Byte(DATAMEM_Byte), 
        .Unsign(DATAMEM_Unsign), .DataOut(MEM_DataOut) );
  RegEn_Nbit32_2 LMDReg ( .A(MEM_DataOut), .Clk(Clk), .Reset(MEMORY_Rst), .EN(
        MEMORY_En), .U(WB_MEM) );
  RegEn_Nbit32_1 WBReg ( .A(MEM_DataIn), .Clk(Clk), .Reset(MEMORY_Rst), .EN(
        MEMORY_En), .U(WB_ALU) );
  RegEn_Nbit5_1 RFWRAddrMEM ( .A(RF_WrAddr_MEM), .Clk(Clk), .Reset(MEMORY_Rst), 
        .EN(MEMORY_En), .U(RF_AddrWR) );
  FD_EN_432 StatusRegMEM ( .D(StatusMEM), .Clk(Clk), .RESET(MEMORY_Rst), .EN(
        MEMORY_En), .Q(\WB_Status[0] ) );
  mux41N_Nbit32_1 WBMux41 ( .in3(WB_MEM), .in2(WB_ALU), .in1({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \WB_Status[0] }), .in0({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .sel(WBMux41_Sel), .Y(RF_DataIn) );
  INV_X1 U3 ( .A(BrZ), .ZN(BrNZ) );
  OR2_X1 U4 ( .A1(Branch_DO), .A2(JRInst_Del), .ZN(FATCHRst_DO) );
endmodule


module DLX ( Clk, Rst );
  input Clk, Rst;
  wire   BrNZ, BrZ, BranchInst, StoreInst, JumpRInst, LHIInst, FATCH_En, Jump,
         DECODE_Rst, DECODE_En, EXECUTE_Rst, EXECUTE_En, MEMORY_Rst, MEMORY_En,
         n1;
  wire   [31:0] Inst;
  wire   [1:0] WBMux41_Sel;
  tri   FS_Rst;
  tri   FATCHRstMux21_Sel;
  tri   [1:0] PCMux41_Sel;
  tri   IRAM_Rst;
  tri   RF_Rst;
  tri   RF_RD1;
  tri   RF_RD2;
  tri   R1Mux21A_Sel;
  tri   R2Mux21B_Sel;
  tri   [1:0] RWMux41WR_Sel;
  tri   ImmMux21_Sel;
  tri   OPAMux21_Sel;
  tri   \OPBMux41_Sel[1] ;
  tri   [3:0] ALU_Sel;
  tri   ALU_Unsign;
  tri   ALU_Arith_logN;
  tri   [2:0] StatusMux81_sel;
  tri   DATAMEM_En;
  tri   DATAMEM_Rst;
  tri   DATAMEM_Read_Wrn;
  tri   DATAMEM_Word;
  tri   DATAMEM_HalfWord;
  tri   DATAMEM_Byte;
  tri   DATAMEM_Unsign;
  tri   RF_WR;
wand  net388923;

  datapath_Nbit32_RAM_DEPTH30_I_SIZE32_DATA_MEM_SIZE10_Nlogicfun3_NALUop4 datap ( 
        .Rst(Rst), .Clk(Clk), .Inst(Inst), .BrNZ(BrNZ), .BrZ(BrZ), 
        .BranchInst(BranchInst), .StoreInst(StoreInst), .JumpRInst(JumpRInst), 
        .LHIInst(LHIInst), .FS_Rst(FS_Rst), .FATCHRstMux21_Sel(
        FATCHRstMux21_Sel), .FATCH_En(FATCH_En), .PCMux41_Sel(PCMux41_Sel), 
        .Jump(Jump), .IRAM_Rst(IRAM_Rst), .DECODE_Rst(DECODE_Rst), .DECODE_En(
        DECODE_En), .RF_Rst(RF_Rst), .RF_RD1(RF_RD1), .RF_RD2(RF_RD2), 
        .R1Mux21A_Sel(R1Mux21A_Sel), .R2Mux21B_Sel(R2Mux21B_Sel), 
        .RWMux41WR_Sel(RWMux41WR_Sel), .ImmMux21_Sel(ImmMux21_Sel), 
        .EXECUTE_Rst(EXECUTE_Rst), .EXECUTE_En(EXECUTE_En), .OPAMux21_Sel(
        OPAMux21_Sel), .OPBMux41_Sel({\OPBMux41_Sel[1] , n1}), .ALU_Sel(
        ALU_Sel), .ALU_Unsign(ALU_Unsign), .ALU_Arith_logN(ALU_Arith_logN), 
        .StatusMux81_sel(StatusMux81_sel), .MEMORY_Rst(MEMORY_Rst), 
        .MEMORY_En(MEMORY_En), .DATAMEM_En(DATAMEM_En), .DATAMEM_Rst(
        DATAMEM_Rst), .DATAMEM_Read_Wrn(DATAMEM_Read_Wrn), .DATAMEM_Word(
        DATAMEM_Word), .DATAMEM_HalfWord(DATAMEM_HalfWord), .DATAMEM_Byte(
        DATAMEM_Byte), .DATAMEM_Unsign(DATAMEM_Unsign), .RF_WR(RF_WR), 
        .WBMux41_Sel(WBMux41_Sel) );
  CU_HW_FUNC_SIZE11_OP_CODE_SIZE6_NALUop4_I_SIZE32_CW_SIZE42 CU ( .Clk(Clk), 
        .Rst(Rst), .Inst(Inst), .BrNZ(BrNZ), .BrZ(BrZ), .BranchInst(BranchInst), .StoreInst(StoreInst), .JumpRInst(JumpRInst), .LHIInst(LHIInst), .FS_Rst(
        FS_Rst), .FATCHRstMux21_Sel(FATCHRstMux21_Sel), .FATCH_En(FATCH_En), 
        .PCMux41_Sel(PCMux41_Sel), .Jump(Jump), .IRAM_Rst(IRAM_Rst), 
        .DECODE_Rst(DECODE_Rst), .DECODE_En(DECODE_En), .RF_Rst(RF_Rst), 
        .RF_RD1(RF_RD1), .RF_RD2(RF_RD2), .R1Mux21A_Sel(R1Mux21A_Sel), 
        .R2Mux21B_Sel(R2Mux21B_Sel), .RWMux41WR_Sel(RWMux41WR_Sel), 
        .ImmMux21_Sel(ImmMux21_Sel), .EXECUTE_Rst(EXECUTE_Rst), .EXECUTE_En(
        EXECUTE_En), .OPAMux21_Sel(OPAMux21_Sel), .OPBMux41_Sel({
        \OPBMux41_Sel[1] , net388923}), .ALU_Sel(ALU_Sel), .ALU_Unsign(
        ALU_Unsign), .ALU_Arith_logN(ALU_Arith_logN), .StatusMux81_sel(
        StatusMux81_sel), .MEMORY_Rst(MEMORY_Rst), .MEMORY_En(MEMORY_En), 
        .DATAMEM_En(DATAMEM_En), .DATAMEM_Rst(DATAMEM_Rst), .DATAMEM_Read_Wrn(
        DATAMEM_Read_Wrn), .DATAMEM_Word(DATAMEM_Word), .DATAMEM_HalfWord(
        DATAMEM_HalfWord), .DATAMEM_Byte(DATAMEM_Byte), .DATAMEM_Unsign(
        DATAMEM_Unsign), .RF_WR(RF_WR), .WBMux41_Sel(WBMux41_Sel) );
  BUF_X2 U1 ( .A(net388923), .Z(n1) );
endmodule

